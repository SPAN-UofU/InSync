// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 10Feb10		Production Release Version 3.1
// SVN Revision Information:
// SVN $Revision: 11146 $
// SVN $Date: 2009-11-21 11:44:53 -0800 (Sat, 21 Nov 2009) $
`timescale 1ns/1ps
module
CoreAHBLite
#
(
parameter
[
5
:
0
]
FAMILY
=
17
,
parameter
[
0
:
0
]
MODE_CFG
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT0ENABLE
=
1
,
parameter
[
0
:
0
]
M0_AHBSLOT1ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT2ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT3ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT4ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT5ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT6ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT7ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT8ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT9ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT10ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT11ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT12ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT13ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT14ENABLE
=
0
,
parameter
[
0
:
0
]
M0_AHBSLOT15ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT0ENABLE
=
1
,
parameter
[
0
:
0
]
M1_AHBSLOT1ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT2ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT3ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT4ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT5ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT6ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT7ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT8ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT9ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT10ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT11ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT12ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT13ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT14ENABLE
=
0
,
parameter
[
0
:
0
]
M1_AHBSLOT15ENABLE
=
0
,
parameter
[
0
:
0
]
M0_HUGESLOTENABLE
=
0
,
parameter
[
0
:
0
]
M1_HUGESLOTENABLE
=
0
,
parameter
[
0
:
0
]
HADDR_SHG_CFG
=
1
,
parameter
[
0
:
0
]
M0_INITCFG0ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG1ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG2ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG3ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG4ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG5ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG6ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG7ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG8ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG9ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG10ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG11ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG12ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG13ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG14ENABLE
=
0
,
parameter
[
0
:
0
]
M0_INITCFG15ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG0ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG1ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG2ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG3ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG4ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG5ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG6ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG7ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG8ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG9ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG10ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG11ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG12ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG13ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG14ENABLE
=
0
,
parameter
[
0
:
0
]
M1_INITCFG15ENABLE
=
0
)
(
input
HCLK,
input
HRESETN,
input
REMAP_M0,
input
[
31
:
0
]
HADDR_M0,
input
HMASTLOCK_M0,
input
[
2
:
0
]
HSIZE_M0,
input
[
1
:
0
]
HTRANS_M0,
input
HWRITE_M0,
input
[
31
:
0
]
HWDATA_M0,
input
[
2
:
0
]
HBURST_M0,
input
[
3
:
0
]
HPROT_M0,
output
wire
[
1
:
0
]
HRESP_M0,
output
wire
[
31
:
0
]
HRDATA_M0,
output
wire
HREADY_M0,
input
[
31
:
0
]
HADDR_M1,
input
HMASTLOCK_M1,
input
[
2
:
0
]
HSIZE_M1,
input
[
1
:
0
]
HTRANS_M1,
input
HWRITE_M1,
input
[
31
:
0
]
HWDATA_M1,
input
[
2
:
0
]
HBURST_M1,
input
[
3
:
0
]
HPROT_M1,
output
wire
[
1
:
0
]
HRESP_M1,
output
wire
[
31
:
0
]
HRDATA_M1,
output
wire
HREADY_M1,
input
[
31
:
0
]
HRDATA_S0,
input
HREADYOUT_S0,
input
[
1
:
0
]
HRESP_S0,
output
wire
HSEL_S0,
output
wire
[
31
:
0
]
HADDR_S0,
output
wire
[
2
:
0
]
HSIZE_S0,
output
wire
[
1
:
0
]
HTRANS_S0,
output
wire
HWRITE_S0,
output
wire
[
31
:
0
]
HWDATA_S0,
output
wire
HREADY_S0,
output
wire
HMASTLOCK_S0,
output
wire
[
2
:
0
]
HBURST_S0,
output
wire
[
3
:
0
]
HPROT_S0,
input
[
31
:
0
]
HRDATA_S1,
input
HREADYOUT_S1,
input
[
1
:
0
]
HRESP_S1,
output
wire
HSEL_S1,
output
wire
[
31
:
0
]
HADDR_S1,
output
wire
[
2
:
0
]
HSIZE_S1,
output
wire
[
1
:
0
]
HTRANS_S1,
output
wire
HWRITE_S1,
output
wire
[
31
:
0
]
HWDATA_S1,
output
wire
HREADY_S1,
output
wire
HMASTLOCK_S1,
output
wire
[
2
:
0
]
HBURST_S1,
output
wire
[
3
:
0
]
HPROT_S1,
input
[
31
:
0
]
HRDATA_S2,
input
HREADYOUT_S2,
input
[
1
:
0
]
HRESP_S2,
output
wire
HSEL_S2,
output
wire
[
31
:
0
]
HADDR_S2,
output
wire
[
2
:
0
]
HSIZE_S2,
output
wire
[
1
:
0
]
HTRANS_S2,
output
wire
HWRITE_S2,
output
wire
[
31
:
0
]
HWDATA_S2,
output
wire
HREADY_S2,
output
wire
HMASTLOCK_S2,
output
wire
[
2
:
0
]
HBURST_S2,
output
wire
[
3
:
0
]
HPROT_S2,
input
[
31
:
0
]
HRDATA_S3,
input
HREADYOUT_S3,
input
[
1
:
0
]
HRESP_S3,
output
wire
HSEL_S3,
output
wire
[
31
:
0
]
HADDR_S3,
output
wire
[
2
:
0
]
HSIZE_S3,
output
wire
[
1
:
0
]
HTRANS_S3,
output
wire
HWRITE_S3,
output
wire
[
31
:
0
]
HWDATA_S3,
output
wire
HREADY_S3,
output
wire
HMASTLOCK_S3,
output
wire
[
2
:
0
]
HBURST_S3,
output
wire
[
3
:
0
]
HPROT_S3,
input
[
31
:
0
]
HRDATA_S4,
input
HREADYOUT_S4,
input
[
1
:
0
]
HRESP_S4,
output
wire
HSEL_S4,
output
wire
[
31
:
0
]
HADDR_S4,
output
wire
[
2
:
0
]
HSIZE_S4,
output
wire
[
1
:
0
]
HTRANS_S4,
output
wire
HWRITE_S4,
output
wire
[
31
:
0
]
HWDATA_S4,
output
wire
HREADY_S4,
output
wire
HMASTLOCK_S4,
output
wire
[
2
:
0
]
HBURST_S4,
output
wire
[
3
:
0
]
HPROT_S4,
input
[
31
:
0
]
HRDATA_S5,
input
HREADYOUT_S5,
input
[
1
:
0
]
HRESP_S5,
output
wire
HSEL_S5,
output
wire
[
31
:
0
]
HADDR_S5,
output
wire
[
2
:
0
]
HSIZE_S5,
output
wire
[
1
:
0
]
HTRANS_S5,
output
wire
HWRITE_S5,
output
wire
[
31
:
0
]
HWDATA_S5,
output
wire
HREADY_S5,
output
wire
HMASTLOCK_S5,
output
wire
[
2
:
0
]
HBURST_S5,
output
wire
[
3
:
0
]
HPROT_S5,
input
[
31
:
0
]
HRDATA_S6,
input
HREADYOUT_S6,
input
[
1
:
0
]
HRESP_S6,
output
wire
HSEL_S6,
output
wire
[
31
:
0
]
HADDR_S6,
output
wire
[
2
:
0
]
HSIZE_S6,
output
wire
[
1
:
0
]
HTRANS_S6,
output
wire
HWRITE_S6,
output
wire
[
31
:
0
]
HWDATA_S6,
output
wire
HREADY_S6,
output
wire
HMASTLOCK_S6,
output
wire
[
2
:
0
]
HBURST_S6,
output
wire
[
3
:
0
]
HPROT_S6,
input
[
31
:
0
]
HRDATA_S7,
input
HREADYOUT_S7,
input
[
1
:
0
]
HRESP_S7,
output
wire
HSEL_S7,
output
wire
[
31
:
0
]
HADDR_S7,
output
wire
[
2
:
0
]
HSIZE_S7,
output
wire
[
1
:
0
]
HTRANS_S7,
output
wire
HWRITE_S7,
output
wire
[
31
:
0
]
HWDATA_S7,
output
wire
HREADY_S7,
output
wire
HMASTLOCK_S7,
output
wire
[
2
:
0
]
HBURST_S7,
output
wire
[
3
:
0
]
HPROT_S7,
input
[
31
:
0
]
HRDATA_S8,
input
HREADYOUT_S8,
input
[
1
:
0
]
HRESP_S8,
output
wire
HSEL_S8,
output
wire
[
31
:
0
]
HADDR_S8,
output
wire
[
2
:
0
]
HSIZE_S8,
output
wire
[
1
:
0
]
HTRANS_S8,
output
wire
HWRITE_S8,
output
wire
[
31
:
0
]
HWDATA_S8,
output
wire
HREADY_S8,
output
wire
HMASTLOCK_S8,
output
wire
[
2
:
0
]
HBURST_S8,
output
wire
[
3
:
0
]
HPROT_S8,
input
[
31
:
0
]
HRDATA_S9,
input
HREADYOUT_S9,
input
[
1
:
0
]
HRESP_S9,
output
wire
HSEL_S9,
output
wire
[
31
:
0
]
HADDR_S9,
output
wire
[
2
:
0
]
HSIZE_S9,
output
wire
[
1
:
0
]
HTRANS_S9,
output
wire
HWRITE_S9,
output
wire
[
31
:
0
]
HWDATA_S9,
output
wire
HREADY_S9,
output
wire
HMASTLOCK_S9,
output
wire
[
2
:
0
]
HBURST_S9,
output
wire
[
3
:
0
]
HPROT_S9,
input
[
31
:
0
]
HRDATA_S10,
input
HREADYOUT_S10,
input
[
1
:
0
]
HRESP_S10,
output
wire
HSEL_S10,
output
wire
[
31
:
0
]
HADDR_S10,
output
wire
[
2
:
0
]
HSIZE_S10,
output
wire
[
1
:
0
]
HTRANS_S10,
output
wire
HWRITE_S10,
output
wire
[
31
:
0
]
HWDATA_S10,
output
wire
HREADY_S10,
output
wire
HMASTLOCK_S10,
output
wire
[
2
:
0
]
HBURST_S10,
output
wire
[
3
:
0
]
HPROT_S10,
input
[
31
:
0
]
HRDATA_S11,
input
HREADYOUT_S11,
input
[
1
:
0
]
HRESP_S11,
output
wire
HSEL_S11,
output
wire
[
31
:
0
]
HADDR_S11,
output
wire
[
2
:
0
]
HSIZE_S11,
output
wire
[
1
:
0
]
HTRANS_S11,
output
wire
HWRITE_S11,
output
wire
[
31
:
0
]
HWDATA_S11,
output
wire
HREADY_S11,
output
wire
HMASTLOCK_S11,
output
wire
[
2
:
0
]
HBURST_S11,
output
wire
[
3
:
0
]
HPROT_S11,
input
[
31
:
0
]
HRDATA_S12,
input
HREADYOUT_S12,
input
[
1
:
0
]
HRESP_S12,
output
wire
HSEL_S12,
output
wire
[
31
:
0
]
HADDR_S12,
output
wire
[
2
:
0
]
HSIZE_S12,
output
wire
[
1
:
0
]
HTRANS_S12,
output
wire
HWRITE_S12,
output
wire
[
31
:
0
]
HWDATA_S12,
output
wire
HREADY_S12,
output
wire
HMASTLOCK_S12,
output
wire
[
2
:
0
]
HBURST_S12,
output
wire
[
3
:
0
]
HPROT_S12,
input
[
31
:
0
]
HRDATA_S13,
input
HREADYOUT_S13,
input
[
1
:
0
]
HRESP_S13,
output
wire
HSEL_S13,
output
wire
[
31
:
0
]
HADDR_S13,
output
wire
[
2
:
0
]
HSIZE_S13,
output
wire
[
1
:
0
]
HTRANS_S13,
output
wire
HWRITE_S13,
output
wire
[
31
:
0
]
HWDATA_S13,
output
wire
HREADY_S13,
output
wire
HMASTLOCK_S13,
output
wire
[
2
:
0
]
HBURST_S13,
output
wire
[
3
:
0
]
HPROT_S13,
input
[
31
:
0
]
HRDATA_S14,
input
HREADYOUT_S14,
input
[
1
:
0
]
HRESP_S14,
output
wire
HSEL_S14,
output
wire
[
31
:
0
]
HADDR_S14,
output
wire
[
2
:
0
]
HSIZE_S14,
output
wire
[
1
:
0
]
HTRANS_S14,
output
wire
HWRITE_S14,
output
wire
[
31
:
0
]
HWDATA_S14,
output
wire
HREADY_S14,
output
wire
HMASTLOCK_S14,
output
wire
[
2
:
0
]
HBURST_S14,
output
wire
[
3
:
0
]
HPROT_S14,
input
[
31
:
0
]
HRDATA_S15,
input
HREADYOUT_S15,
input
[
1
:
0
]
HRESP_S15,
output
wire
HSEL_S15,
output
wire
[
31
:
0
]
HADDR_S15,
output
wire
[
2
:
0
]
HSIZE_S15,
output
wire
[
1
:
0
]
HTRANS_S15,
output
wire
HWRITE_S15,
output
wire
[
31
:
0
]
HWDATA_S15,
output
wire
HREADY_S15,
output
wire
HMASTLOCK_S15,
output
wire
[
2
:
0
]
HBURST_S15,
output
wire
[
3
:
0
]
HPROT_S15,
input
[
31
:
0
]
HRDATA_SHG,
input
HREADYOUT_SHG,
input
[
1
:
0
]
HRESP_SHG,
output
wire
HSEL_SHG,
output
wire
[
31
:
0
]
HADDR_SHG,
output
wire
[
2
:
0
]
HSIZE_SHG,
output
wire
[
1
:
0
]
HTRANS_SHG,
output
wire
HWRITE_SHG,
output
wire
[
31
:
0
]
HWDATA_SHG,
output
wire
HREADY_SHG,
output
wire
HMASTLOCK_SHG,
output
wire
[
2
:
0
]
HBURST_SHG,
output
wire
[
3
:
0
]
HPROT_SHG,
output
wire
INITDATVAL_C0,
output
wire
INITDONE_C0,
output
wire
[
11
:
0
]
INITADDR_C0,
output
wire
[
31
:
0
]
INITDATA_C0,
output
wire
INITDATVAL_C1,
output
wire
INITDONE_C1,
output
wire
[
11
:
0
]
INITADDR_C1,
output
wire
[
31
:
0
]
INITDATA_C1,
output
wire
INITDATVAL_C2,
output
wire
INITDONE_C2,
output
wire
[
11
:
0
]
INITADDR_C2,
output
wire
[
31
:
0
]
INITDATA_C2,
output
wire
INITDATVAL_C3,
output
wire
INITDONE_C3,
output
wire
[
11
:
0
]
INITADDR_C3,
output
wire
[
31
:
0
]
INITDATA_C3,
output
wire
INITDATVAL_C4,
output
wire
INITDONE_C4,
output
wire
[
11
:
0
]
INITADDR_C4,
output
wire
[
31
:
0
]
INITDATA_C4,
output
wire
INITDATVAL_C5,
output
wire
INITDONE_C5,
output
wire
[
11
:
0
]
INITADDR_C5,
output
wire
[
31
:
0
]
INITDATA_C5,
output
wire
INITDATVAL_C6,
output
wire
INITDONE_C6,
output
wire
[
11
:
0
]
INITADDR_C6,
output
wire
[
31
:
0
]
INITDATA_C6,
output
wire
INITDATVAL_C7,
output
wire
INITDONE_C7,
output
wire
[
11
:
0
]
INITADDR_C7,
output
wire
[
31
:
0
]
INITDATA_C7,
output
wire
INITDATVAL_C8,
output
wire
INITDONE_C8,
output
wire
[
11
:
0
]
INITADDR_C8,
output
wire
[
31
:
0
]
INITDATA_C8,
output
wire
INITDATVAL_C9,
output
wire
INITDONE_C9,
output
wire
[
11
:
0
]
INITADDR_C9,
output
wire
[
31
:
0
]
INITDATA_C9,
output
wire
INITDATVAL_C10,
output
wire
INITDONE_C10,
output
wire
[
11
:
0
]
INITADDR_C10,
output
wire
[
31
:
0
]
INITDATA_C10,
output
wire
INITDATVAL_C11,
output
wire
INITDONE_C11,
output
wire
[
11
:
0
]
INITADDR_C11,
output
wire
[
31
:
0
]
INITDATA_C11,
output
wire
INITDATVAL_C12,
output
wire
INITDONE_C12,
output
wire
[
11
:
0
]
INITADDR_C12,
output
wire
[
31
:
0
]
INITDATA_C12,
output
wire
INITDATVAL_C13,
output
wire
INITDONE_C13,
output
wire
[
11
:
0
]
INITADDR_C13,
output
wire
[
31
:
0
]
INITDATA_C13,
output
wire
INITDATVAL_C14,
output
wire
INITDONE_C14,
output
wire
[
11
:
0
]
INITADDR_C14,
output
wire
[
31
:
0
]
INITDATA_C14,
output
wire
INITDATVAL_C15,
output
wire
INITDONE_C15,
output
wire
[
11
:
0
]
INITADDR_C15,
output
wire
[
31
:
0
]
INITDATA_C15
)
;
localparam
[
16
:
0
]
CAHBLTOIl0
=
{
M0_HUGESLOTENABLE
,
M0_AHBSLOT15ENABLE
,
M0_AHBSLOT14ENABLE
,
M0_AHBSLOT13ENABLE
,
M0_AHBSLOT12ENABLE
,
M0_AHBSLOT11ENABLE
,
M0_AHBSLOT10ENABLE
,
M0_AHBSLOT9ENABLE
,
M0_AHBSLOT8ENABLE
,
M0_AHBSLOT7ENABLE
,
M0_AHBSLOT6ENABLE
,
M0_AHBSLOT5ENABLE
,
M0_AHBSLOT4ENABLE
,
M0_AHBSLOT3ENABLE
,
M0_AHBSLOT2ENABLE
,
M0_AHBSLOT1ENABLE
,
M0_AHBSLOT0ENABLE
}
;
localparam
[
16
:
0
]
CAHBLTIIl0
=
{
M1_HUGESLOTENABLE
,
M1_AHBSLOT15ENABLE
,
M1_AHBSLOT14ENABLE
,
M1_AHBSLOT13ENABLE
,
M1_AHBSLOT12ENABLE
,
M1_AHBSLOT11ENABLE
,
M1_AHBSLOT10ENABLE
,
M1_AHBSLOT9ENABLE
,
M1_AHBSLOT8ENABLE
,
M1_AHBSLOT7ENABLE
,
M1_AHBSLOT6ENABLE
,
M1_AHBSLOT5ENABLE
,
M1_AHBSLOT4ENABLE
,
M1_AHBSLOT3ENABLE
,
M1_AHBSLOT2ENABLE
,
M1_AHBSLOT1ENABLE
,
M1_AHBSLOT0ENABLE
}
;
localparam
[
15
:
0
]
CAHBLTO0O0
=
{
M0_INITCFG15ENABLE
,
M0_INITCFG14ENABLE
,
M0_INITCFG13ENABLE
,
M0_INITCFG12ENABLE
,
M0_INITCFG11ENABLE
,
M0_INITCFG10ENABLE
,
M0_INITCFG9ENABLE
,
M0_INITCFG8ENABLE
,
M0_INITCFG7ENABLE
,
M0_INITCFG6ENABLE
,
M0_INITCFG5ENABLE
,
M0_INITCFG4ENABLE
,
M0_INITCFG3ENABLE
,
M0_INITCFG2ENABLE
,
M0_INITCFG1ENABLE
,
M0_INITCFG0ENABLE
}
;
localparam
[
15
:
0
]
CAHBLTI0O0
=
{
M1_INITCFG15ENABLE
,
M1_INITCFG14ENABLE
,
M1_INITCFG13ENABLE
,
M1_INITCFG12ENABLE
,
M1_INITCFG11ENABLE
,
M1_INITCFG10ENABLE
,
M1_INITCFG9ENABLE
,
M1_INITCFG8ENABLE
,
M1_INITCFG7ENABLE
,
M1_INITCFG6ENABLE
,
M1_INITCFG5ENABLE
,
M1_INITCFG4ENABLE
,
M1_INITCFG3ENABLE
,
M1_INITCFG2ENABLE
,
M1_INITCFG1ENABLE
,
M1_INITCFG0ENABLE
}
;
wire
[
31
:
0
]
CAHBLTl0I0l
;
wire
[
15
:
0
]
CAHBLTll0l
;
wire
[
15
:
0
]
CAHBLTO00l
;
wire
[
11
:
0
]
CAHBLTI00l
;
wire
[
31
:
0
]
CAHBLTl00l
;
assign
HTRANS_S0
[
0
]
=
1
'b
0
;
assign
HTRANS_S1
[
0
]
=
1
'b
0
;
assign
HTRANS_S2
[
0
]
=
1
'b
0
;
assign
HTRANS_S3
[
0
]
=
1
'b
0
;
assign
HTRANS_S4
[
0
]
=
1
'b
0
;
assign
HTRANS_S5
[
0
]
=
1
'b
0
;
assign
HTRANS_S6
[
0
]
=
1
'b
0
;
assign
HTRANS_S7
[
0
]
=
1
'b
0
;
assign
HTRANS_S8
[
0
]
=
1
'b
0
;
assign
HTRANS_S9
[
0
]
=
1
'b
0
;
assign
HTRANS_S10
[
0
]
=
1
'b
0
;
assign
HTRANS_S11
[
0
]
=
1
'b
0
;
assign
HTRANS_S12
[
0
]
=
1
'b
0
;
assign
HTRANS_S13
[
0
]
=
1
'b
0
;
assign
HTRANS_S14
[
0
]
=
1
'b
0
;
assign
HTRANS_S15
[
0
]
=
1
'b
0
;
assign
HTRANS_SHG
[
0
]
=
1
'b
0
;
assign
HRESP_M0
[
1
]
=
1
'b
0
;
assign
HRESP_M1
[
1
]
=
1
'b
0
;
assign
HBURST_S0
=
3
'b
0
;
assign
HBURST_S1
=
3
'b
0
;
assign
HBURST_S2
=
3
'b
0
;
assign
HBURST_S3
=
3
'b
0
;
assign
HBURST_S4
=
3
'b
0
;
assign
HBURST_S5
=
3
'b
0
;
assign
HBURST_S6
=
3
'b
0
;
assign
HBURST_S7
=
3
'b
0
;
assign
HBURST_S8
=
3
'b
0
;
assign
HBURST_S9
=
3
'b
0
;
assign
HBURST_S10
=
3
'b
0
;
assign
HBURST_S11
=
3
'b
0
;
assign
HBURST_S12
=
3
'b
0
;
assign
HBURST_S13
=
3
'b
0
;
assign
HBURST_S14
=
3
'b
0
;
assign
HBURST_S15
=
3
'b
0
;
assign
HBURST_SHG
=
3
'b
0
;
assign
HPROT_S0
=
4
'b
0
;
assign
HPROT_S1
=
4
'b
0
;
assign
HPROT_S2
=
4
'b
0
;
assign
HPROT_S3
=
4
'b
0
;
assign
HPROT_S4
=
4
'b
0
;
assign
HPROT_S5
=
4
'b
0
;
assign
HPROT_S6
=
4
'b
0
;
assign
HPROT_S7
=
4
'b
0
;
assign
HPROT_S8
=
4
'b
0
;
assign
HPROT_S9
=
4
'b
0
;
assign
HPROT_S10
=
4
'b
0
;
assign
HPROT_S11
=
4
'b
0
;
assign
HPROT_S12
=
4
'b
0
;
assign
HPROT_S13
=
4
'b
0
;
assign
HPROT_S14
=
4
'b
0
;
assign
HPROT_S15
=
4
'b
0
;
assign
HPROT_SHG
=
4
'b
0
;
CAHBLTlOl0
#
(
.MODE_CFG
(
MODE_CFG
)
,
.CAHBLTOIl0
(
CAHBLTOIl0
)
,
.CAHBLTIIl0
(
CAHBLTIIl0
)
,
.CAHBLTO0O0
(
CAHBLTO0O0
)
,
.CAHBLTI0O0
(
CAHBLTI0O0
)
)
CAHBLTO1I0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.REMAP_M0
(
REMAP_M0
)
,
.HADDR_M0
(
HADDR_M0
)
,
.HMASTLOCK_M0
(
HMASTLOCK_M0
)
,
.HSIZE_M0
(
HSIZE_M0
)
,
.HTRANS_M0
(
HTRANS_M0
[
1
]
)
,
.HWRITE_M0
(
HWRITE_M0
)
,
.HWDATA_M0
(
HWDATA_M0
)
,
.HRESP_M0
(
HRESP_M0
[
0
]
)
,
.HRDATA_M0
(
HRDATA_M0
)
,
.HREADY_M0
(
HREADY_M0
)
,
.HADDR_M1
(
HADDR_M1
)
,
.HMASTLOCK_M1
(
HMASTLOCK_M1
)
,
.HSIZE_M1
(
HSIZE_M1
)
,
.HTRANS_M1
(
HTRANS_M1
[
1
]
)
,
.HWRITE_M1
(
HWRITE_M1
)
,
.HWDATA_M1
(
HWDATA_M1
)
,
.HRESP_M1
(
HRESP_M1
[
0
]
)
,
.HRDATA_M1
(
HRDATA_M1
)
,
.HREADY_M1
(
HREADY_M1
)
,
.HRDATA_S0
(
HRDATA_S0
)
,
.HREADYOUT_S0
(
HREADYOUT_S0
)
,
.HRESP_S0
(
HRESP_S0
[
0
]
)
,
.HSEL_S0
(
HSEL_S0
)
,
.HADDR_S0
(
HADDR_S0
)
,
.HSIZE_S0
(
HSIZE_S0
)
,
.HTRANS_S0
(
HTRANS_S0
[
1
]
)
,
.HWRITE_S0
(
HWRITE_S0
)
,
.HWDATA_S0
(
HWDATA_S0
)
,
.HREADY_S0
(
HREADY_S0
)
,
.HMASTLOCK_S0
(
HMASTLOCK_S0
)
,
.HRDATA_S1
(
HRDATA_S1
)
,
.HREADYOUT_S1
(
HREADYOUT_S1
)
,
.HRESP_S1
(
HRESP_S1
[
0
]
)
,
.HSEL_S1
(
HSEL_S1
)
,
.HADDR_S1
(
HADDR_S1
)
,
.HSIZE_S1
(
HSIZE_S1
)
,
.HTRANS_S1
(
HTRANS_S1
[
1
]
)
,
.HWRITE_S1
(
HWRITE_S1
)
,
.HWDATA_S1
(
HWDATA_S1
)
,
.HREADY_S1
(
HREADY_S1
)
,
.HMASTLOCK_S1
(
HMASTLOCK_S1
)
,
.HRDATA_S2
(
HRDATA_S2
)
,
.HREADYOUT_S2
(
HREADYOUT_S2
)
,
.HRESP_S2
(
HRESP_S2
[
0
]
)
,
.HSEL_S2
(
HSEL_S2
)
,
.HADDR_S2
(
HADDR_S2
)
,
.HSIZE_S2
(
HSIZE_S2
)
,
.HTRANS_S2
(
HTRANS_S2
[
1
]
)
,
.HWRITE_S2
(
HWRITE_S2
)
,
.HWDATA_S2
(
HWDATA_S2
)
,
.HREADY_S2
(
HREADY_S2
)
,
.HMASTLOCK_S2
(
HMASTLOCK_S2
)
,
.HRDATA_S3
(
HRDATA_S3
)
,
.HREADYOUT_S3
(
HREADYOUT_S3
)
,
.HRESP_S3
(
HRESP_S3
[
0
]
)
,
.HSEL_S3
(
HSEL_S3
)
,
.HADDR_S3
(
HADDR_S3
)
,
.HSIZE_S3
(
HSIZE_S3
)
,
.HTRANS_S3
(
HTRANS_S3
[
1
]
)
,
.HWRITE_S3
(
HWRITE_S3
)
,
.HWDATA_S3
(
HWDATA_S3
)
,
.HREADY_S3
(
HREADY_S3
)
,
.HMASTLOCK_S3
(
HMASTLOCK_S3
)
,
.HRDATA_S4
(
HRDATA_S4
)
,
.HREADYOUT_S4
(
HREADYOUT_S4
)
,
.HRESP_S4
(
HRESP_S4
[
0
]
)
,
.HSEL_S4
(
HSEL_S4
)
,
.HADDR_S4
(
HADDR_S4
)
,
.HSIZE_S4
(
HSIZE_S4
)
,
.HTRANS_S4
(
HTRANS_S4
[
1
]
)
,
.HWRITE_S4
(
HWRITE_S4
)
,
.HWDATA_S4
(
HWDATA_S4
)
,
.HREADY_S4
(
HREADY_S4
)
,
.HMASTLOCK_S4
(
HMASTLOCK_S4
)
,
.HRDATA_S5
(
HRDATA_S5
)
,
.HREADYOUT_S5
(
HREADYOUT_S5
)
,
.HRESP_S5
(
HRESP_S5
[
0
]
)
,
.HSEL_S5
(
HSEL_S5
)
,
.HADDR_S5
(
HADDR_S5
)
,
.HSIZE_S5
(
HSIZE_S5
)
,
.HTRANS_S5
(
HTRANS_S5
[
1
]
)
,
.HWRITE_S5
(
HWRITE_S5
)
,
.HWDATA_S5
(
HWDATA_S5
)
,
.HREADY_S5
(
HREADY_S5
)
,
.HMASTLOCK_S5
(
HMASTLOCK_S5
)
,
.HRDATA_S6
(
HRDATA_S6
)
,
.HREADYOUT_S6
(
HREADYOUT_S6
)
,
.HRESP_S6
(
HRESP_S6
[
0
]
)
,
.HSEL_S6
(
HSEL_S6
)
,
.HADDR_S6
(
HADDR_S6
)
,
.HSIZE_S6
(
HSIZE_S6
)
,
.HTRANS_S6
(
HTRANS_S6
[
1
]
)
,
.HWRITE_S6
(
HWRITE_S6
)
,
.HWDATA_S6
(
HWDATA_S6
)
,
.HREADY_S6
(
HREADY_S6
)
,
.HMASTLOCK_S6
(
HMASTLOCK_S6
)
,
.HRDATA_S7
(
HRDATA_S7
)
,
.HREADYOUT_S7
(
HREADYOUT_S7
)
,
.HRESP_S7
(
HRESP_S7
[
0
]
)
,
.HSEL_S7
(
HSEL_S7
)
,
.HADDR_S7
(
HADDR_S7
)
,
.HSIZE_S7
(
HSIZE_S7
)
,
.HTRANS_S7
(
HTRANS_S7
[
1
]
)
,
.HWRITE_S7
(
HWRITE_S7
)
,
.HWDATA_S7
(
HWDATA_S7
)
,
.HREADY_S7
(
HREADY_S7
)
,
.HMASTLOCK_S7
(
HMASTLOCK_S7
)
,
.HRDATA_S8
(
HRDATA_S8
)
,
.HREADYOUT_S8
(
HREADYOUT_S8
)
,
.HRESP_S8
(
HRESP_S8
[
0
]
)
,
.HSEL_S8
(
HSEL_S8
)
,
.HADDR_S8
(
HADDR_S8
)
,
.HSIZE_S8
(
HSIZE_S8
)
,
.HTRANS_S8
(
HTRANS_S8
[
1
]
)
,
.HWRITE_S8
(
HWRITE_S8
)
,
.HWDATA_S8
(
HWDATA_S8
)
,
.HREADY_S8
(
HREADY_S8
)
,
.HMASTLOCK_S8
(
HMASTLOCK_S8
)
,
.HRDATA_S9
(
HRDATA_S9
)
,
.HREADYOUT_S9
(
HREADYOUT_S9
)
,
.HRESP_S9
(
HRESP_S9
[
0
]
)
,
.HSEL_S9
(
HSEL_S9
)
,
.HADDR_S9
(
HADDR_S9
)
,
.HSIZE_S9
(
HSIZE_S9
)
,
.HTRANS_S9
(
HTRANS_S9
[
1
]
)
,
.HWRITE_S9
(
HWRITE_S9
)
,
.HWDATA_S9
(
HWDATA_S9
)
,
.HREADY_S9
(
HREADY_S9
)
,
.HMASTLOCK_S9
(
HMASTLOCK_S9
)
,
.HRDATA_S10
(
HRDATA_S10
)
,
.HREADYOUT_S10
(
HREADYOUT_S10
)
,
.HRESP_S10
(
HRESP_S10
[
0
]
)
,
.HSEL_S10
(
HSEL_S10
)
,
.HADDR_S10
(
HADDR_S10
)
,
.HSIZE_S10
(
HSIZE_S10
)
,
.HTRANS_S10
(
HTRANS_S10
[
1
]
)
,
.HWRITE_S10
(
HWRITE_S10
)
,
.HWDATA_S10
(
HWDATA_S10
)
,
.HREADY_S10
(
HREADY_S10
)
,
.HMASTLOCK_S10
(
HMASTLOCK_S10
)
,
.HRDATA_S11
(
HRDATA_S11
)
,
.HREADYOUT_S11
(
HREADYOUT_S11
)
,
.HRESP_S11
(
HRESP_S11
[
0
]
)
,
.HSEL_S11
(
HSEL_S11
)
,
.HADDR_S11
(
HADDR_S11
)
,
.HSIZE_S11
(
HSIZE_S11
)
,
.HTRANS_S11
(
HTRANS_S11
[
1
]
)
,
.HWRITE_S11
(
HWRITE_S11
)
,
.HWDATA_S11
(
HWDATA_S11
)
,
.HREADY_S11
(
HREADY_S11
)
,
.HMASTLOCK_S11
(
HMASTLOCK_S11
)
,
.HRDATA_S12
(
HRDATA_S12
)
,
.HREADYOUT_S12
(
HREADYOUT_S12
)
,
.HRESP_S12
(
HRESP_S12
[
0
]
)
,
.HSEL_S12
(
HSEL_S12
)
,
.HADDR_S12
(
HADDR_S12
)
,
.HSIZE_S12
(
HSIZE_S12
)
,
.HTRANS_S12
(
HTRANS_S12
[
1
]
)
,
.HWRITE_S12
(
HWRITE_S12
)
,
.HWDATA_S12
(
HWDATA_S12
)
,
.HREADY_S12
(
HREADY_S12
)
,
.HMASTLOCK_S12
(
HMASTLOCK_S12
)
,
.HRDATA_S13
(
HRDATA_S13
)
,
.HREADYOUT_S13
(
HREADYOUT_S13
)
,
.HRESP_S13
(
HRESP_S13
[
0
]
)
,
.HSEL_S13
(
HSEL_S13
)
,
.HADDR_S13
(
HADDR_S13
)
,
.HSIZE_S13
(
HSIZE_S13
)
,
.HTRANS_S13
(
HTRANS_S13
[
1
]
)
,
.HWRITE_S13
(
HWRITE_S13
)
,
.HWDATA_S13
(
HWDATA_S13
)
,
.HREADY_S13
(
HREADY_S13
)
,
.HMASTLOCK_S13
(
HMASTLOCK_S13
)
,
.HRDATA_S14
(
HRDATA_S14
)
,
.HREADYOUT_S14
(
HREADYOUT_S14
)
,
.HRESP_S14
(
HRESP_S14
[
0
]
)
,
.HSEL_S14
(
HSEL_S14
)
,
.HADDR_S14
(
HADDR_S14
)
,
.HSIZE_S14
(
HSIZE_S14
)
,
.HTRANS_S14
(
HTRANS_S14
[
1
]
)
,
.HWRITE_S14
(
HWRITE_S14
)
,
.HWDATA_S14
(
HWDATA_S14
)
,
.HREADY_S14
(
HREADY_S14
)
,
.HMASTLOCK_S14
(
HMASTLOCK_S14
)
,
.HRDATA_S15
(
HRDATA_S15
)
,
.HREADYOUT_S15
(
HREADYOUT_S15
)
,
.HRESP_S15
(
HRESP_S15
[
0
]
)
,
.HSEL_S15
(
HSEL_S15
)
,
.HADDR_S15
(
HADDR_S15
)
,
.HSIZE_S15
(
HSIZE_S15
)
,
.HTRANS_S15
(
HTRANS_S15
[
1
]
)
,
.HWRITE_S15
(
HWRITE_S15
)
,
.HWDATA_S15
(
HWDATA_S15
)
,
.HREADY_S15
(
HREADY_S15
)
,
.HMASTLOCK_S15
(
HMASTLOCK_S15
)
,
.HRDATA_SHG
(
HRDATA_SHG
)
,
.HREADYOUT_SHG
(
HREADYOUT_SHG
)
,
.HRESP_SHG
(
HRESP_SHG
[
0
]
)
,
.HSEL_SHG
(
HSEL_SHG
)
,
.HADDR_SHG
(
CAHBLTl0I0l
)
,
.HSIZE_SHG
(
HSIZE_SHG
)
,
.HTRANS_SHG
(
HTRANS_SHG
[
1
]
)
,
.HWRITE_SHG
(
HWRITE_SHG
)
,
.HWDATA_SHG
(
HWDATA_SHG
)
,
.HREADY_SHG
(
HREADY_SHG
)
,
.HMASTLOCK_SHG
(
HMASTLOCK_SHG
)
,
.CAHBLTll0l
(
CAHBLTll0l
)
,
.CAHBLTO00l
(
CAHBLTO00l
)
,
.CAHBLTI00l
(
CAHBLTI00l
)
,
.CAHBLTl00l
(
CAHBLTl00l
)
)
;
assign
{
INITDATVAL_C15
,
INITDATVAL_C14
,
INITDATVAL_C13
,
INITDATVAL_C12
,
INITDATVAL_C11
,
INITDATVAL_C10
,
INITDATVAL_C9
,
INITDATVAL_C8
,
INITDATVAL_C7
,
INITDATVAL_C6
,
INITDATVAL_C5
,
INITDATVAL_C4
,
INITDATVAL_C3
,
INITDATVAL_C2
,
INITDATVAL_C1
,
INITDATVAL_C0
}
=
CAHBLTll0l
[
15
:
0
]
;
assign
{
INITDONE_C15
,
INITDONE_C14
,
INITDONE_C13
,
INITDONE_C12
,
INITDONE_C11
,
INITDONE_C10
,
INITDONE_C9
,
INITDONE_C8
,
INITDONE_C7
,
INITDONE_C6
,
INITDONE_C5
,
INITDONE_C4
,
INITDONE_C3
,
INITDONE_C2
,
INITDONE_C1
,
INITDONE_C0
}
=
CAHBLTO00l
[
15
:
0
]
;
assign
{
INITADDR_C15
[
11
:
0
]
,
INITADDR_C14
[
11
:
0
]
,
INITADDR_C13
[
11
:
0
]
,
INITADDR_C12
[
11
:
0
]
,
INITADDR_C11
[
11
:
0
]
,
INITADDR_C10
[
11
:
0
]
,
INITADDR_C9
[
11
:
0
]
,
INITADDR_C8
[
11
:
0
]
,
INITADDR_C7
[
11
:
0
]
,
INITADDR_C6
[
11
:
0
]
,
INITADDR_C5
[
11
:
0
]
,
INITADDR_C4
[
11
:
0
]
,
INITADDR_C3
[
11
:
0
]
,
INITADDR_C2
[
11
:
0
]
,
INITADDR_C1
[
11
:
0
]
,
INITADDR_C0
[
11
:
0
]
}
=
{
16
{
CAHBLTI00l
[
11
:
0
]
}
}
;
assign
{
INITDATA_C15
[
31
:
0
]
,
INITDATA_C14
[
31
:
0
]
,
INITDATA_C13
[
31
:
0
]
,
INITDATA_C12
[
31
:
0
]
,
INITDATA_C11
[
31
:
0
]
,
INITDATA_C10
[
31
:
0
]
,
INITDATA_C9
[
31
:
0
]
,
INITDATA_C8
[
31
:
0
]
,
INITDATA_C7
[
31
:
0
]
,
INITDATA_C6
[
31
:
0
]
,
INITDATA_C5
[
31
:
0
]
,
INITDATA_C4
[
31
:
0
]
,
INITDATA_C3
[
31
:
0
]
,
INITDATA_C2
[
31
:
0
]
,
INITDATA_C1
[
31
:
0
]
,
INITDATA_C0
[
31
:
0
]
}
=
{
16
{
CAHBLTl00l
[
31
:
0
]
}
}
;
generate
begin
:
CAHBLTI1I0l
if
(
MODE_CFG
==
0
)
begin
:
CAHBLTlI0
assign
HADDR_SHG
[
31
]
=
CAHBLTl0I0l
[
31
]
;
end
else
if
(
MODE_CFG
==
1
)
begin
:
CAHBLTIl0
if
(
HADDR_SHG_CFG
==
0
)
begin
:
CAHBLTl1I0l
assign
HADDR_SHG
[
31
]
=
1
'b
0
;
end
else
if
(
HADDR_SHG_CFG
==
1
)
begin
:
CAHBLTOOl0l
assign
HADDR_SHG
[
31
]
=
1
'b
1
;
end
end
end
endgenerate
assign
HADDR_SHG
[
30
:
0
]
=
CAHBLTl0I0l
[
30
:
0
]
;
endmodule
