// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 10Feb10		Production Release Version 3.1
// SVN Revision Information:
// SVN $Revision: 11955 $
// SVN $Date: 2010-01-30 15:35:13 -0800 (Sat, 30 Jan 2010) $
`timescale 1ns/1ps
module
CAHBLTlOl0
#
(
parameter
[
0
:
0
]
MODE_CFG
=
0
,
parameter
[
16
:
0
]
CAHBLTOIl0
=
(
2
**
17
)
-
1
,
parameter
[
16
:
0
]
CAHBLTIIl0
=
(
2
**
17
)
-
1
,
parameter
[
15
:
0
]
CAHBLTO0O0
=
0
,
parameter
[
15
:
0
]
CAHBLTI0O0
=
0
)
(
input
HCLK,
input
HRESETN,
input
REMAP_M0,
input
[
31
:
0
]
HADDR_M0,
input
HMASTLOCK_M0,
input
[
2
:
0
]
HSIZE_M0,
input
HTRANS_M0,
input
HWRITE_M0,
input
[
31
:
0
]
HWDATA_M0,
output
wire
HRESP_M0,
output
wire
[
31
:
0
]
HRDATA_M0,
output
wire
HREADY_M0,
input
[
31
:
0
]
HADDR_M1,
input
HMASTLOCK_M1,
input
[
2
:
0
]
HSIZE_M1,
input
HTRANS_M1,
input
HWRITE_M1,
input
[
31
:
0
]
HWDATA_M1,
output
wire
HRESP_M1,
output
wire
[
31
:
0
]
HRDATA_M1,
output
wire
HREADY_M1,
input
[
31
:
0
]
HRDATA_S0,
input
HREADYOUT_S0,
input
HRESP_S0,
output
wire
HSEL_S0,
output
wire
[
31
:
0
]
HADDR_S0,
output
wire
[
2
:
0
]
HSIZE_S0,
output
wire
HTRANS_S0,
output
wire
HWRITE_S0,
output
wire
[
31
:
0
]
HWDATA_S0,
output
wire
HREADY_S0,
output
wire
HMASTLOCK_S0,
input
[
31
:
0
]
HRDATA_S1,
input
HREADYOUT_S1,
input
HRESP_S1,
output
wire
HSEL_S1,
output
wire
[
31
:
0
]
HADDR_S1,
output
wire
[
2
:
0
]
HSIZE_S1,
output
wire
HTRANS_S1,
output
wire
HWRITE_S1,
output
wire
[
31
:
0
]
HWDATA_S1,
output
wire
HREADY_S1,
output
wire
HMASTLOCK_S1,
input
[
31
:
0
]
HRDATA_S2,
input
HREADYOUT_S2,
input
HRESP_S2,
output
wire
HSEL_S2,
output
wire
[
31
:
0
]
HADDR_S2,
output
wire
[
2
:
0
]
HSIZE_S2,
output
wire
HTRANS_S2,
output
wire
HWRITE_S2,
output
wire
[
31
:
0
]
HWDATA_S2,
output
wire
HREADY_S2,
output
wire
HMASTLOCK_S2,
input
[
31
:
0
]
HRDATA_S3,
input
HREADYOUT_S3,
input
HRESP_S3,
output
wire
HSEL_S3,
output
wire
[
31
:
0
]
HADDR_S3,
output
wire
[
2
:
0
]
HSIZE_S3,
output
wire
HTRANS_S3,
output
wire
HWRITE_S3,
output
wire
[
31
:
0
]
HWDATA_S3,
output
wire
HREADY_S3,
output
wire
HMASTLOCK_S3,
input
[
31
:
0
]
HRDATA_S4,
input
HREADYOUT_S4,
input
HRESP_S4,
output
wire
HSEL_S4,
output
wire
[
31
:
0
]
HADDR_S4,
output
wire
[
2
:
0
]
HSIZE_S4,
output
wire
HTRANS_S4,
output
wire
HWRITE_S4,
output
wire
[
31
:
0
]
HWDATA_S4,
output
wire
HREADY_S4,
output
wire
HMASTLOCK_S4,
input
[
31
:
0
]
HRDATA_S5,
input
HREADYOUT_S5,
input
HRESP_S5,
output
wire
HSEL_S5,
output
wire
[
31
:
0
]
HADDR_S5,
output
wire
[
2
:
0
]
HSIZE_S5,
output
wire
HTRANS_S5,
output
wire
HWRITE_S5,
output
wire
[
31
:
0
]
HWDATA_S5,
output
wire
HREADY_S5,
output
wire
HMASTLOCK_S5,
input
[
31
:
0
]
HRDATA_S6,
input
HREADYOUT_S6,
input
HRESP_S6,
output
wire
HSEL_S6,
output
wire
[
31
:
0
]
HADDR_S6,
output
wire
[
2
:
0
]
HSIZE_S6,
output
wire
HTRANS_S6,
output
wire
HWRITE_S6,
output
wire
[
31
:
0
]
HWDATA_S6,
output
wire
HREADY_S6,
output
wire
HMASTLOCK_S6,
input
[
31
:
0
]
HRDATA_S7,
input
HREADYOUT_S7,
input
HRESP_S7,
output
wire
HSEL_S7,
output
wire
[
31
:
0
]
HADDR_S7,
output
wire
[
2
:
0
]
HSIZE_S7,
output
wire
HTRANS_S7,
output
wire
HWRITE_S7,
output
wire
[
31
:
0
]
HWDATA_S7,
output
wire
HREADY_S7,
output
wire
HMASTLOCK_S7,
input
[
31
:
0
]
HRDATA_S8,
input
HREADYOUT_S8,
input
HRESP_S8,
output
wire
HSEL_S8,
output
wire
[
31
:
0
]
HADDR_S8,
output
wire
[
2
:
0
]
HSIZE_S8,
output
wire
HTRANS_S8,
output
wire
HWRITE_S8,
output
wire
[
31
:
0
]
HWDATA_S8,
output
wire
HREADY_S8,
output
wire
HMASTLOCK_S8,
input
[
31
:
0
]
HRDATA_S9,
input
HREADYOUT_S9,
input
HRESP_S9,
output
wire
HSEL_S9,
output
wire
[
31
:
0
]
HADDR_S9,
output
wire
[
2
:
0
]
HSIZE_S9,
output
wire
HTRANS_S9,
output
wire
HWRITE_S9,
output
wire
[
31
:
0
]
HWDATA_S9,
output
wire
HREADY_S9,
output
wire
HMASTLOCK_S9,
input
[
31
:
0
]
HRDATA_S10,
input
HREADYOUT_S10,
input
HRESP_S10,
output
wire
HSEL_S10,
output
wire
[
31
:
0
]
HADDR_S10,
output
wire
[
2
:
0
]
HSIZE_S10,
output
wire
HTRANS_S10,
output
wire
HWRITE_S10,
output
wire
[
31
:
0
]
HWDATA_S10,
output
wire
HREADY_S10,
output
wire
HMASTLOCK_S10,
input
[
31
:
0
]
HRDATA_S11,
input
HREADYOUT_S11,
input
HRESP_S11,
output
wire
HSEL_S11,
output
wire
[
31
:
0
]
HADDR_S11,
output
wire
[
2
:
0
]
HSIZE_S11,
output
wire
HTRANS_S11,
output
wire
HWRITE_S11,
output
wire
[
31
:
0
]
HWDATA_S11,
output
wire
HREADY_S11,
output
wire
HMASTLOCK_S11,
input
[
31
:
0
]
HRDATA_S12,
input
HREADYOUT_S12,
input
HRESP_S12,
output
wire
HSEL_S12,
output
wire
[
31
:
0
]
HADDR_S12,
output
wire
[
2
:
0
]
HSIZE_S12,
output
wire
HTRANS_S12,
output
wire
HWRITE_S12,
output
wire
[
31
:
0
]
HWDATA_S12,
output
wire
HREADY_S12,
output
wire
HMASTLOCK_S12,
input
[
31
:
0
]
HRDATA_S13,
input
HREADYOUT_S13,
input
HRESP_S13,
output
wire
HSEL_S13,
output
wire
[
31
:
0
]
HADDR_S13,
output
wire
[
2
:
0
]
HSIZE_S13,
output
wire
HTRANS_S13,
output
wire
HWRITE_S13,
output
wire
[
31
:
0
]
HWDATA_S13,
output
wire
HREADY_S13,
output
wire
HMASTLOCK_S13,
input
[
31
:
0
]
HRDATA_S14,
input
HREADYOUT_S14,
input
HRESP_S14,
output
wire
HSEL_S14,
output
wire
[
31
:
0
]
HADDR_S14,
output
wire
[
2
:
0
]
HSIZE_S14,
output
wire
HTRANS_S14,
output
wire
HWRITE_S14,
output
wire
[
31
:
0
]
HWDATA_S14,
output
wire
HREADY_S14,
output
wire
HMASTLOCK_S14,
input
[
31
:
0
]
HRDATA_S15,
input
HREADYOUT_S15,
input
HRESP_S15,
output
wire
HSEL_S15,
output
wire
[
31
:
0
]
HADDR_S15,
output
wire
[
2
:
0
]
HSIZE_S15,
output
wire
HTRANS_S15,
output
wire
HWRITE_S15,
output
wire
[
31
:
0
]
HWDATA_S15,
output
wire
HREADY_S15,
output
wire
HMASTLOCK_S15,
input
[
31
:
0
]
HRDATA_SHG,
input
HREADYOUT_SHG,
input
HRESP_SHG,
output
wire
HSEL_SHG,
output
wire
[
31
:
0
]
HADDR_SHG,
output
wire
[
2
:
0
]
HSIZE_SHG,
output
wire
HTRANS_SHG,
output
wire
HWRITE_SHG,
output
wire
[
31
:
0
]
HWDATA_SHG,
output
wire
HREADY_SHG,
output
wire
HMASTLOCK_SHG,
output
wire
[
15
:
0
]
CAHBLTll0l,
output
wire
[
15
:
0
]
CAHBLTO00l,
output
wire
[
11
:
0
]
CAHBLTI00l,
output
wire
[
31
:
0
]
CAHBLTl00l
)
;
wire
[
31
:
0
]
CAHBLTOlll
;
wire
CAHBLTll1
;
wire
[
2
:
0
]
CAHBLTIlll
;
wire
CAHBLTllll
;
wire
CAHBLTO0ll
;
wire
CAHBLTlIl0
;
wire
CAHBLTOll0
;
wire
CAHBLTIll0
;
wire
CAHBLTlll0
;
wire
CAHBLTO0l0
;
wire
CAHBLTI0l0
;
wire
CAHBLTl0l0
;
wire
CAHBLTO1l0
;
wire
CAHBLTI1l0
;
wire
CAHBLTl1l0
;
wire
CAHBLTOO00
;
wire
CAHBLTIO00
;
wire
CAHBLTlO00
;
wire
CAHBLTOI00
;
wire
CAHBLTII00
;
wire
CAHBLTlI00
;
wire
CAHBLTOl00
;
wire
CAHBLTIl00
;
wire
CAHBLTll00
;
wire
CAHBLTO000
;
wire
CAHBLTI000
;
wire
CAHBLTl000
;
wire
CAHBLTO100
;
wire
CAHBLTI100
;
wire
CAHBLTl100
;
wire
CAHBLTOO10
;
wire
CAHBLTIO10
;
wire
CAHBLTlO10
;
wire
CAHBLTOI10
;
wire
CAHBLTII10
;
wire
CAHBLTlI10
;
wire
CAHBLTOl10
;
wire
CAHBLTIl10
;
wire
CAHBLTll10
;
wire
CAHBLTO010
;
wire
CAHBLTI010
;
wire
CAHBLTl010
;
wire
CAHBLTO110
;
wire
CAHBLTI110
;
wire
CAHBLTl110
;
wire
CAHBLTOOO1
;
wire
CAHBLTIOO1
;
wire
CAHBLTlOO1
;
wire
CAHBLTOIO1
;
wire
CAHBLTIIO1
;
wire
CAHBLTlIO1
;
wire
CAHBLTOlO1
;
wire
CAHBLTIlO1
;
wire
CAHBLTllO1
;
wire
CAHBLTO0O1
;
wire
CAHBLTI0O1
;
wire
CAHBLTl0O1
;
wire
CAHBLTO1O1
;
wire
CAHBLTI1O1
;
wire
CAHBLTl1O1
;
wire
CAHBLTOOI1
;
wire
CAHBLTIOI1
;
wire
CAHBLTlOI1
;
wire
CAHBLTOII1
;
wire
CAHBLTIII1
;
wire
CAHBLTlII1
;
wire
CAHBLTOlI1
;
wire
CAHBLTIlI1
;
wire
CAHBLTllI1
;
wire
CAHBLTO0I1
;
wire
CAHBLTI0I1
;
wire
CAHBLTl0I1
;
wire
CAHBLTO1I1
;
wire
CAHBLTI1I1
;
wire
CAHBLTl1I1
;
wire
CAHBLTOOl1
;
wire
CAHBLTIOl1
;
wire
CAHBLTlOl1
;
wire
CAHBLTOIl1
;
wire
CAHBLTIIl1
;
wire
CAHBLTlIl1
;
wire
CAHBLTOll1
;
wire
CAHBLTIll1
;
wire
CAHBLTlll1
;
wire
CAHBLTO0l1
;
wire
CAHBLTI0l1
;
wire
CAHBLTl0l1
;
wire
CAHBLTO1l1
;
wire
CAHBLTI1l1
;
wire
CAHBLTl1l1
;
wire
CAHBLTOO01
;
wire
CAHBLTIO01
;
wire
CAHBLTlO01
;
wire
CAHBLTOI01
;
wire
CAHBLTII01
;
wire
CAHBLTlI01
;
wire
CAHBLTOl01
;
wire
CAHBLTIl01
;
wire
CAHBLTll01
;
wire
CAHBLTO001
;
wire
CAHBLTI001
;
wire
CAHBLTl001
;
wire
CAHBLTO101
;
wire
CAHBLTI101
;
wire
CAHBLTl101
;
wire
CAHBLTOO11
;
wire
CAHBLTIO11
;
wire
CAHBLTlO11
;
wire
CAHBLTOI11
;
wire
CAHBLTII11
;
wire
CAHBLTlI11
;
wire
CAHBLTOl11
;
wire
CAHBLTIl11
;
wire
CAHBLTll11
;
wire
CAHBLTO011
;
wire
CAHBLTI011
;
wire
CAHBLTl011
;
wire
CAHBLTO111
;
wire
CAHBLTI111
;
wire
CAHBLTl111
;
wire
CAHBLTOOOOI
;
wire
CAHBLTIOOOI
;
wire
CAHBLTlOOOI
;
wire
CAHBLTOIOOI
;
wire
CAHBLTIIOOI
;
wire
CAHBLTlIOOI
;
wire
CAHBLTOlOOI
;
wire
CAHBLTIlOOI
;
wire
CAHBLTllOOI
;
wire
CAHBLTO0OOI
;
wire
CAHBLTI0OOI
;
wire
CAHBLTl0OOI
;
wire
CAHBLTO1OOI
;
wire
CAHBLTI1OOI
;
wire
CAHBLTl1OOI
;
wire
CAHBLTOOIOI
;
wire
CAHBLTIOIOI
;
wire
CAHBLTlOIOI
;
wire
CAHBLTOIIOI
;
wire
CAHBLTIIIOI
;
wire
CAHBLTlIIOI
;
wire
CAHBLTOlIOI
;
wire
CAHBLTIlIOI
;
wire
CAHBLTllIOI
;
wire
CAHBLTO0IOI
;
wire
CAHBLTI0IOI
;
wire
CAHBLTl0IOI
;
wire
CAHBLTO1IOI
;
wire
CAHBLTI1IOI
;
wire
CAHBLTl1IOI
;
wire
CAHBLTOOlOI
;
wire
CAHBLTIOlOI
;
wire
CAHBLTlOlOI
;
wire
CAHBLTOIlOI
;
wire
CAHBLTIIlOI
;
wire
CAHBLTlIlOI
;
wire
CAHBLTOllOI
;
wire
CAHBLTIllOI
;
wire
CAHBLTlllOI
;
wire
CAHBLTO0lOI
;
wire
CAHBLTI0lOI
;
wire
CAHBLTl0lOI
;
wire
CAHBLTO1lOI
;
wire
CAHBLTI1lOI
;
wire
CAHBLTl1lOI
;
wire
CAHBLTOO0OI
;
wire
CAHBLTIO0OI
;
wire
CAHBLTlO0OI
;
wire
CAHBLTOI0OI
;
wire
CAHBLTII0OI
;
wire
CAHBLTlI0OI
;
wire
CAHBLTOl0OI
;
wire
CAHBLTIl0OI
;
wire
CAHBLTll0OI
;
wire
CAHBLTO00OI
;
wire
CAHBLTI00OI
;
wire
CAHBLTl00OI
;
wire
CAHBLTO10OI
;
wire
CAHBLTI10OI
;
wire
CAHBLTl10OI
;
wire
CAHBLTOO1OI
;
wire
CAHBLTIO1OI
;
wire
CAHBLTlO1OI
;
wire
CAHBLTOI1OI
;
wire
CAHBLTII1OI
;
wire
CAHBLTlI1OI
;
wire
[
31
:
0
]
CAHBLTI0ll
;
wire
CAHBLTO01
;
wire
[
2
:
0
]
CAHBLTl0ll
;
wire
CAHBLTO1ll
;
wire
CAHBLTI1ll
;
wire
CAHBLTOl1OI
;
wire
CAHBLTIl1OI
;
wire
CAHBLTll1OI
;
wire
CAHBLTO01OI
;
wire
CAHBLTI01OI
;
wire
CAHBLTl01OI
;
wire
CAHBLTO11OI
;
wire
CAHBLTI11OI
;
wire
CAHBLTl11OI
;
wire
CAHBLTOOOII
;
wire
CAHBLTIOOII
;
wire
CAHBLTlOOII
;
wire
CAHBLTOIOII
;
wire
CAHBLTIIOII
;
wire
CAHBLTlIOII
;
wire
CAHBLTOlOII
;
wire
CAHBLTIlOII
;
wire
CAHBLTllOII
;
wire
CAHBLTO0OII
;
wire
CAHBLTI0OII
;
wire
CAHBLTl0OII
;
wire
CAHBLTO1OII
;
wire
CAHBLTI1OII
;
wire
CAHBLTl1OII
;
wire
CAHBLTOOIII
;
wire
CAHBLTIOIII
;
wire
CAHBLTlOIII
;
wire
CAHBLTOIIII
;
wire
CAHBLTIIIII
;
wire
CAHBLTlIIII
;
wire
CAHBLTOlIII
;
wire
CAHBLTIlIII
;
wire
CAHBLTllIII
;
wire
CAHBLTO0III
;
wire
CAHBLTI0III
;
wire
CAHBLTl0III
;
wire
CAHBLTO1III
;
wire
CAHBLTI1III
;
wire
CAHBLTl1III
;
wire
CAHBLTOOlII
;
wire
CAHBLTIOlII
;
wire
CAHBLTlOlII
;
wire
CAHBLTOIlII
;
wire
CAHBLTIIlII
;
wire
CAHBLTlIlII
;
wire
CAHBLTOllII
;
wire
CAHBLTIllII
;
wire
CAHBLTlllII
;
wire
CAHBLTO0lII
;
wire
CAHBLTI0lII
;
wire
CAHBLTl0lII
;
wire
CAHBLTO1lII
;
wire
CAHBLTI1lII
;
wire
CAHBLTl1lII
;
wire
CAHBLTOO0II
;
wire
CAHBLTIO0II
;
wire
CAHBLTlO0II
;
wire
CAHBLTOI0II
;
wire
CAHBLTII0II
;
wire
CAHBLTlI0II
;
wire
CAHBLTOl0II
;
wire
CAHBLTIl0II
;
wire
CAHBLTll0II
;
wire
CAHBLTO00II
;
wire
CAHBLTI00II
;
wire
CAHBLTl00II
;
wire
CAHBLTO10II
;
wire
CAHBLTI10II
;
wire
CAHBLTl10II
;
wire
CAHBLTOO1II
;
wire
CAHBLTIO1II
;
wire
CAHBLTlO1II
;
wire
CAHBLTOI1II
;
wire
CAHBLTII1II
;
wire
CAHBLTlI1II
;
wire
CAHBLTOl1II
;
wire
CAHBLTIl1II
;
wire
CAHBLTll1II
;
wire
CAHBLTO01II
;
wire
CAHBLTI01II
;
wire
CAHBLTl01II
;
wire
CAHBLTO11II
;
wire
CAHBLTI11II
;
wire
CAHBLTl11II
;
wire
CAHBLTOOOlI
;
wire
CAHBLTIOOlI
;
wire
CAHBLTlOOlI
;
wire
CAHBLTOIOlI
;
wire
CAHBLTIIOlI
;
wire
CAHBLTlIOlI
;
wire
CAHBLTOlOlI
;
wire
CAHBLTIlOlI
;
wire
CAHBLTllOlI
;
wire
CAHBLTO0OlI
;
wire
CAHBLTI0OlI
;
wire
CAHBLTl0OlI
;
wire
CAHBLTO1OlI
;
wire
CAHBLTI1OlI
;
wire
CAHBLTl1OlI
;
wire
CAHBLTOOIlI
;
wire
CAHBLTIOIlI
;
wire
CAHBLTlOIlI
;
wire
CAHBLTOIIlI
;
wire
CAHBLTIIIlI
;
wire
CAHBLTlIIlI
;
wire
CAHBLTOlIlI
;
wire
CAHBLTIlIlI
;
wire
CAHBLTllIlI
;
wire
CAHBLTO0IlI
;
wire
CAHBLTI0IlI
;
wire
CAHBLTl0IlI
;
wire
CAHBLTO1IlI
;
wire
CAHBLTI1IlI
;
wire
CAHBLTl1IlI
;
wire
CAHBLTOOllI
;
wire
CAHBLTIOllI
;
wire
CAHBLTlOllI
;
wire
CAHBLTOIllI
;
wire
CAHBLTIIllI
;
wire
CAHBLTlIllI
;
wire
CAHBLTOlllI
;
wire
CAHBLTIlllI
;
wire
CAHBLTllllI
;
wire
CAHBLTO0llI
;
wire
CAHBLTI0llI
;
wire
CAHBLTl0llI
;
wire
CAHBLTO1llI
;
wire
CAHBLTI1llI
;
wire
CAHBLTl1llI
;
wire
CAHBLTOO0lI
;
wire
CAHBLTIO0lI
;
wire
CAHBLTlO0lI
;
wire
CAHBLTOI0lI
;
wire
CAHBLTII0lI
;
wire
CAHBLTlI0lI
;
wire
CAHBLTOl0lI
;
wire
CAHBLTIl0lI
;
wire
CAHBLTll0lI
;
wire
CAHBLTO00lI
;
wire
CAHBLTI00lI
;
wire
CAHBLTl00lI
;
wire
CAHBLTO10lI
;
wire
CAHBLTI10lI
;
wire
CAHBLTl10lI
;
wire
CAHBLTOO1lI
;
wire
CAHBLTIO1lI
;
wire
CAHBLTlO1lI
;
wire
CAHBLTOI1lI
;
wire
CAHBLTII1lI
;
wire
CAHBLTlI1lI
;
wire
CAHBLTOl1lI
;
wire
CAHBLTIl1lI
;
wire
CAHBLTll1lI
;
wire
CAHBLTO01lI
;
wire
CAHBLTI01lI
;
wire
CAHBLTl01lI
;
wire
CAHBLTO11lI
;
wire
CAHBLTI11lI
;
wire
CAHBLTl11lI
;
wire
CAHBLTOOO0I
;
wire
CAHBLTIOO0I
;
wire
CAHBLTlOO0I
;
wire
CAHBLTOIO0I
;
wire
CAHBLTIIO0I
;
wire
CAHBLTlIO0I
;
wire
CAHBLTOlO0I
;
wire
CAHBLTIlO0I
;
wire
CAHBLTllO0I
;
wire
CAHBLTO0O0I
;
wire
CAHBLTI0O0I
;
wire
CAHBLTl0O0I
;
wire
CAHBLTO1O0I
;
wire
CAHBLTI1O0I
;
wire
CAHBLTl1O0I
;
wire
CAHBLTOOI0I
;
wire
CAHBLTIOI0I
;
wire
CAHBLTlOI0I
;
wire
CAHBLTOII0I
;
wire
CAHBLTIII0I
;
wire
CAHBLTlII0I
;
wire
CAHBLTOlI0I
;
wire
CAHBLTIlI0I
;
wire
[
15
:
0
]
CAHBLTl0O0
;
wire
[
15
:
0
]
CAHBLTO1O0
;
wire
[
31
:
0
]
CAHBLTllI0I
;
wire
[
31
:
0
]
CAHBLTO0I0I
;
wire
[
31
:
0
]
CAHBLTI0I0I
;
wire
[
31
:
0
]
CAHBLTl0I0I
;
wire
[
31
:
0
]
CAHBLTO1I0I
;
wire
[
31
:
0
]
CAHBLTI1I0I
;
wire
[
31
:
0
]
CAHBLTl1I0I
;
wire
[
31
:
0
]
CAHBLTOOl0I
;
wire
[
31
:
0
]
CAHBLTIOl0I
;
wire
[
31
:
0
]
CAHBLTlOl0I
;
wire
[
31
:
0
]
CAHBLTOIl0I
;
wire
[
31
:
0
]
CAHBLTIIl0I
;
wire
[
31
:
0
]
CAHBLTlIl0I
;
wire
[
31
:
0
]
CAHBLTOll0I
;
wire
[
31
:
0
]
CAHBLTIll0I
;
wire
[
31
:
0
]
CAHBLTlll0I
;
wire
[
31
:
0
]
CAHBLTO0l0I
;
wire
[
31
:
0
]
CAHBLTI0l0I
;
wire
[
31
:
0
]
CAHBLTl0l0I
;
wire
[
31
:
0
]
CAHBLTO1l0I
;
wire
[
31
:
0
]
CAHBLTI1l0I
;
wire
[
31
:
0
]
CAHBLTl1l0I
;
wire
[
31
:
0
]
CAHBLTOO00I
;
wire
[
31
:
0
]
CAHBLTIO00I
;
wire
[
31
:
0
]
CAHBLTlO00I
;
wire
[
31
:
0
]
CAHBLTOI00I
;
wire
[
31
:
0
]
CAHBLTII00I
;
wire
[
31
:
0
]
CAHBLTlI00I
;
wire
[
31
:
0
]
CAHBLTOl00I
;
wire
[
31
:
0
]
CAHBLTIl00I
;
wire
[
31
:
0
]
CAHBLTll00I
;
wire
[
31
:
0
]
CAHBLTO000I
;
wire
[
31
:
0
]
CAHBLTI000I
;
wire
[
31
:
0
]
CAHBLTl000I
;
wire
CAHBLTO100I
;
wire
CAHBLTI100I
;
wire
CAHBLTl100I
;
wire
CAHBLTOO10I
;
wire
CAHBLTIO10I
;
wire
CAHBLTlO10I
;
wire
CAHBLTOI10I
;
wire
CAHBLTII10I
;
wire
CAHBLTlI10I
;
wire
CAHBLTOl10I
;
wire
CAHBLTIl10I
;
wire
CAHBLTll10I
;
wire
CAHBLTO010I
;
wire
CAHBLTI010I
;
wire
CAHBLTl010I
;
wire
CAHBLTO110I
;
wire
CAHBLTI110I
;
wire
CAHBLTl110I
;
wire
CAHBLTOOO1I
;
wire
CAHBLTIOO1I
;
wire
CAHBLTlOO1I
;
wire
CAHBLTOIO1I
;
wire
CAHBLTIIO1I
;
wire
CAHBLTlIO1I
;
wire
CAHBLTOlO1I
;
wire
CAHBLTIlO1I
;
wire
CAHBLTllO1I
;
wire
CAHBLTO0O1I
;
wire
CAHBLTI0O1I
;
wire
CAHBLTl0O1I
;
wire
CAHBLTO1O1I
;
wire
CAHBLTI1O1I
;
wire
CAHBLTl1O1I
;
wire
CAHBLTOOI1I
;
wire
CAHBLTIOI1I
;
wire
CAHBLTlOI1I
;
wire
CAHBLTOII1I
;
wire
CAHBLTIII1I
;
wire
CAHBLTlII1I
;
wire
CAHBLTOlI1I
;
wire
CAHBLTIlI1I
;
wire
CAHBLTllI1I
;
wire
CAHBLTO0I1I
;
wire
CAHBLTI0I1I
;
wire
CAHBLTl0I1I
;
wire
CAHBLTO1I1I
;
wire
CAHBLTI1I1I
;
wire
CAHBLTl1I1I
;
wire
CAHBLTOOl1I
;
wire
CAHBLTIOl1I
;
wire
CAHBLTlOl1I
;
wire
CAHBLTOIl1I
;
wire
CAHBLTIIl1I
;
wire
CAHBLTlIl1I
;
wire
CAHBLTOll1I
;
wire
CAHBLTIll1I
;
wire
CAHBLTlll1I
;
wire
CAHBLTO0l1I
;
wire
CAHBLTI0l1I
;
wire
CAHBLTl0l1I
;
wire
CAHBLTO1l1I
;
wire
CAHBLTI1l1I
;
wire
CAHBLTl1l1I
;
wire
CAHBLTOO01I
;
wire
CAHBLTIO01I
;
wire
CAHBLTlO01I
;
wire
CAHBLTOI01I
;
wire
CAHBLTII01I
;
wire
CAHBLTlI01I
;
wire
CAHBLTOl01I
;
wire
[
31
:
0
]
CAHBLTIl01I
;
wire
[
31
:
0
]
CAHBLTll01I
;
wire
[
31
:
0
]
CAHBLTO001I
;
wire
[
31
:
0
]
CAHBLTI001I
;
wire
[
31
:
0
]
CAHBLTl001I
;
wire
[
31
:
0
]
CAHBLTO101I
;
wire
[
31
:
0
]
CAHBLTI101I
;
wire
[
31
:
0
]
CAHBLTl101I
;
wire
[
31
:
0
]
CAHBLTOO11I
;
wire
[
31
:
0
]
CAHBLTIO11I
;
wire
[
31
:
0
]
CAHBLTlO11I
;
wire
[
31
:
0
]
CAHBLTOI11I
;
wire
[
31
:
0
]
CAHBLTII11I
;
wire
[
31
:
0
]
CAHBLTlI11I
;
wire
[
31
:
0
]
CAHBLTOl11I
;
wire
[
31
:
0
]
CAHBLTIl11I
;
wire
[
31
:
0
]
CAHBLTll11I
;
wire
[
31
:
0
]
CAHBLTO011I
;
wire
[
31
:
0
]
CAHBLTI011I
;
wire
[
31
:
0
]
CAHBLTl011I
;
wire
[
31
:
0
]
CAHBLTO111I
;
wire
[
31
:
0
]
CAHBLTI111I
;
wire
[
31
:
0
]
CAHBLTl111I
;
wire
[
31
:
0
]
CAHBLTOOOOl
;
wire
[
31
:
0
]
CAHBLTIOOOl
;
wire
[
31
:
0
]
CAHBLTlOOOl
;
wire
[
31
:
0
]
CAHBLTOIOOl
;
wire
[
31
:
0
]
CAHBLTIIOOl
;
wire
[
31
:
0
]
CAHBLTlIOOl
;
wire
[
31
:
0
]
CAHBLTOlOOl
;
wire
[
31
:
0
]
CAHBLTIlOOl
;
wire
[
31
:
0
]
CAHBLTllOOl
;
wire
[
31
:
0
]
CAHBLTO0OOl
;
wire
[
31
:
0
]
CAHBLTI0OOl
;
wire
[
31
:
0
]
CAHBLTl0OOl
;
wire
[
31
:
0
]
CAHBLTO1OOl
;
wire
[
31
:
0
]
CAHBLTI1OOl
;
wire
[
31
:
0
]
CAHBLTl1OOl
;
wire
[
31
:
0
]
CAHBLTOOIOl
;
wire
[
31
:
0
]
CAHBLTIOIOl
;
wire
[
31
:
0
]
CAHBLTlOIOl
;
wire
[
31
:
0
]
CAHBLTOIIOl
;
wire
[
31
:
0
]
CAHBLTIIIOl
;
wire
[
31
:
0
]
CAHBLTlIIOl
;
wire
[
31
:
0
]
CAHBLTOlIOl
;
wire
[
31
:
0
]
CAHBLTIlIOl
;
wire
[
31
:
0
]
CAHBLTllIOl
;
wire
[
31
:
0
]
CAHBLTO0IOl
;
wire
[
31
:
0
]
CAHBLTI0IOl
;
wire
[
31
:
0
]
CAHBLTl0IOl
;
wire
[
31
:
0
]
CAHBLTO1IOl
;
wire
[
31
:
0
]
CAHBLTI1IOl
;
wire
[
31
:
0
]
CAHBLTl1IOl
;
wire
[
31
:
0
]
CAHBLTOOlOl
;
wire
[
31
:
0
]
CAHBLTIOlOl
;
wire
[
31
:
0
]
CAHBLTlOlOl
;
wire
[
31
:
0
]
CAHBLTOIlOl
;
wire
[
31
:
0
]
CAHBLTIIlOl
;
wire
[
31
:
0
]
CAHBLTlIlOl
;
wire
[
31
:
0
]
CAHBLTOllOl
;
wire
[
31
:
0
]
CAHBLTIllOl
;
wire
[
31
:
0
]
CAHBLTlllOl
;
wire
[
31
:
0
]
CAHBLTO0lOl
;
wire
[
31
:
0
]
CAHBLTI0lOl
;
wire
[
31
:
0
]
CAHBLTl0lOl
;
wire
[
31
:
0
]
CAHBLTO1lOl
;
wire
[
31
:
0
]
CAHBLTI1lOl
;
wire
[
31
:
0
]
CAHBLTl1lOl
;
wire
[
31
:
0
]
CAHBLTOO0Ol
;
wire
[
31
:
0
]
CAHBLTIO0Ol
;
wire
[
31
:
0
]
CAHBLTlO0Ol
;
wire
[
31
:
0
]
CAHBLTOI0Ol
;
wire
[
2
:
0
]
CAHBLTII0Ol
;
wire
[
2
:
0
]
CAHBLTlI0Ol
;
wire
[
2
:
0
]
CAHBLTOl0Ol
;
wire
[
2
:
0
]
CAHBLTIl0Ol
;
wire
[
2
:
0
]
CAHBLTll0Ol
;
wire
[
2
:
0
]
CAHBLTO00Ol
;
wire
[
2
:
0
]
CAHBLTI00Ol
;
wire
[
2
:
0
]
CAHBLTl00Ol
;
wire
[
2
:
0
]
CAHBLTO10Ol
;
wire
[
2
:
0
]
CAHBLTI10Ol
;
wire
[
2
:
0
]
CAHBLTl10Ol
;
wire
[
2
:
0
]
CAHBLTOO1Ol
;
wire
[
2
:
0
]
CAHBLTIO1Ol
;
wire
[
2
:
0
]
CAHBLTlO1Ol
;
wire
[
2
:
0
]
CAHBLTOI1Ol
;
wire
[
2
:
0
]
CAHBLTII1Ol
;
wire
[
2
:
0
]
CAHBLTlI1Ol
;
wire
[
2
:
0
]
CAHBLTOl1Ol
;
wire
[
2
:
0
]
CAHBLTIl1Ol
;
wire
[
2
:
0
]
CAHBLTll1Ol
;
wire
[
2
:
0
]
CAHBLTO01Ol
;
wire
[
2
:
0
]
CAHBLTI01Ol
;
wire
[
2
:
0
]
CAHBLTl01Ol
;
wire
[
2
:
0
]
CAHBLTO11Ol
;
wire
[
2
:
0
]
CAHBLTI11Ol
;
wire
[
2
:
0
]
CAHBLTl11Ol
;
wire
[
2
:
0
]
CAHBLTOOOIl
;
wire
[
2
:
0
]
CAHBLTIOOIl
;
wire
[
2
:
0
]
CAHBLTlOOIl
;
wire
[
2
:
0
]
CAHBLTOIOIl
;
wire
[
2
:
0
]
CAHBLTIIOIl
;
wire
[
2
:
0
]
CAHBLTlIOIl
;
wire
[
2
:
0
]
CAHBLTOlOIl
;
wire
[
2
:
0
]
CAHBLTIlOIl
;
wire
[
2
:
0
]
CAHBLTllOIl
;
wire
[
2
:
0
]
CAHBLTO0OIl
;
wire
CAHBLTI0OIl
;
wire
CAHBLTl0OIl
;
wire
CAHBLTO1OIl
;
wire
CAHBLTI1OIl
;
wire
CAHBLTl1OIl
;
wire
CAHBLTOOIIl
;
wire
CAHBLTIOIIl
;
wire
CAHBLTlOIIl
;
wire
CAHBLTOIIIl
;
wire
CAHBLTIIIIl
;
wire
CAHBLTlIIIl
;
wire
CAHBLTOlIIl
;
wire
CAHBLTIlIIl
;
wire
CAHBLTllIIl
;
wire
CAHBLTO0IIl
;
wire
CAHBLTI0IIl
;
wire
CAHBLTl0IIl
;
wire
CAHBLTO1IIl
;
wire
CAHBLTI1IIl
;
wire
CAHBLTl1IIl
;
wire
CAHBLTOOlIl
;
wire
CAHBLTIOlIl
;
wire
CAHBLTlOlIl
;
wire
CAHBLTOIlIl
;
wire
CAHBLTIIlIl
;
wire
CAHBLTlIlIl
;
wire
CAHBLTOllIl
;
wire
CAHBLTIllIl
;
wire
CAHBLTlllIl
;
wire
CAHBLTO0lIl
;
wire
CAHBLTI0lIl
;
wire
CAHBLTl0lIl
;
wire
CAHBLTO1lIl
;
wire
CAHBLTI1lIl
;
wire
CAHBLTl1lIl
;
wire
CAHBLTOO0Il
;
wire
CAHBLTIO0Il
;
wire
CAHBLTlO0Il
;
wire
CAHBLTOI0Il
;
wire
CAHBLTII0Il
;
wire
CAHBLTlI0Il
;
wire
CAHBLTOl0Il
;
wire
CAHBLTIl0Il
;
wire
CAHBLTll0Il
;
wire
CAHBLTO00Il
;
wire
CAHBLTI00Il
;
wire
CAHBLTl00Il
;
wire
CAHBLTO10Il
;
wire
CAHBLTI10Il
;
wire
CAHBLTl10Il
;
wire
CAHBLTOO1Il
;
wire
CAHBLTIO1Il
;
wire
CAHBLTlO1Il
;
wire
CAHBLTOI1Il
;
wire
CAHBLTII1Il
;
wire
CAHBLTlI1Il
;
wire
CAHBLTOl1Il
;
wire
CAHBLTIl1Il
;
wire
CAHBLTll1Il
;
wire
CAHBLTO01Il
;
wire
CAHBLTI01Il
;
wire
CAHBLTl01Il
;
wire
CAHBLTO11Il
;
wire
CAHBLTI11Il
;
wire
CAHBLTl11Il
;
wire
CAHBLTOOOll
;
wire
CAHBLTIOOll
;
wire
CAHBLTlOOll
;
wire
CAHBLTOIOll
;
wire
CAHBLTIIOll
;
wire
CAHBLTlIOll
;
wire
CAHBLTOlOll
;
wire
CAHBLTIlOll
;
wire
CAHBLTllOll
;
wire
CAHBLTO0Oll
;
wire
CAHBLTI0Oll
;
wire
CAHBLTl0Oll
;
wire
CAHBLTO1Oll
;
wire
CAHBLTI1Oll
;
wire
CAHBLTl1Oll
;
wire
CAHBLTOOIll
;
wire
CAHBLTIOIll
;
wire
CAHBLTlOIll
;
wire
CAHBLTOIIll
;
wire
CAHBLTIIIll
;
wire
CAHBLTlIIll
;
wire
CAHBLTOlIll
;
wire
CAHBLTIlIll
;
wire
CAHBLTllIll
;
wire
CAHBLTO0Ill
;
wire
CAHBLTI0Ill
;
wire
CAHBLTl0Ill
;
wire
CAHBLTO1Ill
;
wire
CAHBLTI1Ill
;
wire
CAHBLTl1Ill
;
wire
CAHBLTOOlll
;
wire
CAHBLTIOlll
;
wire
CAHBLTlOlll
;
wire
CAHBLTOIlll
;
wire
CAHBLTIIlll
;
wire
CAHBLTlIlll
;
wire
CAHBLTOllll
;
wire
CAHBLTIllll
;
wire
CAHBLTlllll
;
wire
CAHBLTO0lll
;
wire
CAHBLTI0lll
;
wire
CAHBLTl0lll
;
wire
CAHBLTO1lll
;
wire
CAHBLTI1lll
;
wire
CAHBLTl1lll
;
wire
CAHBLTOO0ll
;
wire
CAHBLTIO0ll
;
wire
CAHBLTlO0ll
;
wire
CAHBLTOI0ll
;
wire
CAHBLTII0ll
;
wire
CAHBLTlI0ll
;
wire
CAHBLTOl0ll
;
wire
CAHBLTIl0ll
;
wire
CAHBLTll0ll
;
wire
CAHBLTO00ll
;
wire
CAHBLTI00ll
;
wire
CAHBLTl00ll
;
wire
CAHBLTO10ll
;
wire
CAHBLTI10ll
;
wire
CAHBLTl10ll
;
wire
CAHBLTOO1ll
;
wire
CAHBLTIO1ll
;
wire
CAHBLTlO1ll
;
wire
CAHBLTOI1ll
;
wire
CAHBLTII1ll
;
wire
CAHBLTlI1ll
;
wire
CAHBLTOl1ll
;
wire
CAHBLTIl1ll
;
wire
CAHBLTll1ll
;
wire
CAHBLTO01ll
;
wire
CAHBLTI01ll
;
wire
CAHBLTl01ll
;
wire
CAHBLTO11ll
;
wire
CAHBLTI11ll
;
wire
CAHBLTl11ll
;
wire
CAHBLTOOO0l
;
wire
CAHBLTIOO0l
;
wire
CAHBLTlOO0l
;
wire
CAHBLTOIO0l
;
wire
CAHBLTIIO0l
;
wire
CAHBLTlIO0l
;
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTI1l0
=
CAHBLTlll0
;
else
assign
CAHBLTI1l0
=
1
'b
1
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTll00
=
CAHBLTOI00
;
else
assign
CAHBLTll00
=
1
'b
1
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTOI10
=
CAHBLTI100
;
else
assign
CAHBLTOI10
=
1
'b
1
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTI110
=
CAHBLTll10
;
else
assign
CAHBLTI110
=
1
'b
1
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTllO1
=
CAHBLTOIO1
;
else
assign
CAHBLTllO1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTOII1
=
CAHBLTI1O1
;
else
assign
CAHBLTOII1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTI1I1
=
CAHBLTllI1
;
else
assign
CAHBLTI1I1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTlll1
=
CAHBLTOIl1
;
else
assign
CAHBLTlll1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTOI01
=
CAHBLTI1l1
;
else
assign
CAHBLTOI01
=
1
'b
1
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTI101
=
CAHBLTll01
;
else
assign
CAHBLTI101
=
1
'b
1
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTll11
=
CAHBLTOI11
;
else
assign
CAHBLTll11
=
1
'b
1
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTOIOOI
=
CAHBLTI111
;
else
assign
CAHBLTOIOOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTI1OOI
=
CAHBLTllOOI
;
else
assign
CAHBLTI1OOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTllIOI
=
CAHBLTOIIOI
;
else
assign
CAHBLTllIOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTOIlOI
=
CAHBLTI1IOI
;
else
assign
CAHBLTOIlOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTI1lOI
=
CAHBLTlllOI
;
else
assign
CAHBLTI1lOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTll0OI
=
CAHBLTOI0OI
;
else
assign
CAHBLTll0OI
=
1
'b
1
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOI1OI
=
CAHBLTI10OI
;
else
assign
CAHBLTOI1OI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTl11OI
=
CAHBLTO01OI
;
else
assign
CAHBLTl11OI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTO0OII
=
CAHBLTIIOII
;
else
assign
CAHBLTO0OII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTIIIII
=
CAHBLTl1OII
;
else
assign
CAHBLTIIIII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTl1III
=
CAHBLTO0III
;
else
assign
CAHBLTl1III
=
1
'b
1
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTO0lII
=
CAHBLTIIlII
;
else
assign
CAHBLTO0lII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTII0II
=
CAHBLTl1lII
;
else
assign
CAHBLTII0II
=
1
'b
1
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTl10II
=
CAHBLTO00II
;
else
assign
CAHBLTl10II
=
1
'b
1
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTO01II
=
CAHBLTII1II
;
else
assign
CAHBLTO01II
=
1
'b
1
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTIIOlI
=
CAHBLTl11II
;
else
assign
CAHBLTIIOlI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTl1OlI
=
CAHBLTO0OlI
;
else
assign
CAHBLTl1OlI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTO0IlI
=
CAHBLTIIIlI
;
else
assign
CAHBLTO0IlI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTIIllI
=
CAHBLTl1IlI
;
else
assign
CAHBLTIIllI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTl1llI
=
CAHBLTO0llI
;
else
assign
CAHBLTl1llI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTO00lI
=
CAHBLTII0lI
;
else
assign
CAHBLTO00lI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTII1lI
=
CAHBLTl10lI
;
else
assign
CAHBLTII1lI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTl11lI
=
CAHBLTO01lI
;
else
assign
CAHBLTl11lI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTO0O0I
=
CAHBLTIIO0I
;
else
assign
CAHBLTO0O0I
=
1
'b
1
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTIII0I
=
CAHBLTl1O0I
;
else
assign
CAHBLTIII0I
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTl1l0
=
CAHBLTO0l0
;
else
assign
CAHBLTl1l0
=
1
'b
1
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTO000
=
CAHBLTII00
;
else
assign
CAHBLTO000
=
1
'b
1
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTII10
=
CAHBLTl100
;
else
assign
CAHBLTII10
=
1
'b
1
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTl110
=
CAHBLTO010
;
else
assign
CAHBLTl110
=
1
'b
1
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTO0O1
=
CAHBLTIIO1
;
else
assign
CAHBLTO0O1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTIII1
=
CAHBLTl1O1
;
else
assign
CAHBLTIII1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTl1I1
=
CAHBLTO0I1
;
else
assign
CAHBLTl1I1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTO0l1
=
CAHBLTIIl1
;
else
assign
CAHBLTO0l1
=
1
'b
1
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTII01
=
CAHBLTl1l1
;
else
assign
CAHBLTII01
=
1
'b
1
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTl101
=
CAHBLTO001
;
else
assign
CAHBLTl101
=
1
'b
1
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTO011
=
CAHBLTII11
;
else
assign
CAHBLTO011
=
1
'b
1
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTIIOOI
=
CAHBLTl111
;
else
assign
CAHBLTIIOOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTl1OOI
=
CAHBLTO0OOI
;
else
assign
CAHBLTl1OOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTO0IOI
=
CAHBLTIIIOI
;
else
assign
CAHBLTO0IOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTIIlOI
=
CAHBLTl1IOI
;
else
assign
CAHBLTIIlOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTl1lOI
=
CAHBLTO0lOI
;
else
assign
CAHBLTl1lOI
=
1
'b
1
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTO00OI
=
CAHBLTII0OI
;
else
assign
CAHBLTO00OI
=
1
'b
1
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTII1OI
=
CAHBLTl10OI
;
else
assign
CAHBLTII1OI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTOOOII
=
CAHBLTI01OI
;
else
assign
CAHBLTOOOII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTI0OII
=
CAHBLTlIOII
;
else
assign
CAHBLTI0OII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTlIIII
=
CAHBLTOOIII
;
else
assign
CAHBLTlIIII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTOOlII
=
CAHBLTI0III
;
else
assign
CAHBLTOOlII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTI0lII
=
CAHBLTlIlII
;
else
assign
CAHBLTI0lII
=
1
'b
1
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTlI0II
=
CAHBLTOO0II
;
else
assign
CAHBLTlI0II
=
1
'b
1
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTOO1II
=
CAHBLTI00II
;
else
assign
CAHBLTOO1II
=
1
'b
1
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTI01II
=
CAHBLTlI1II
;
else
assign
CAHBLTI01II
=
1
'b
1
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTlIOlI
=
CAHBLTOOOlI
;
else
assign
CAHBLTlIOlI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTOOIlI
=
CAHBLTI0OlI
;
else
assign
CAHBLTOOIlI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTI0IlI
=
CAHBLTlIIlI
;
else
assign
CAHBLTI0IlI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTlIllI
=
CAHBLTOOllI
;
else
assign
CAHBLTlIllI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTOO0lI
=
CAHBLTI0llI
;
else
assign
CAHBLTOO0lI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTI00lI
=
CAHBLTlI0lI
;
else
assign
CAHBLTI00lI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTlI1lI
=
CAHBLTOO1lI
;
else
assign
CAHBLTlI1lI
=
1
'b
1
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTOOO0I
=
CAHBLTI01lI
;
else
assign
CAHBLTOOO0I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTI0O0I
=
CAHBLTlIO0I
;
else
assign
CAHBLTI0O0I
=
1
'b
1
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTlII0I
=
CAHBLTOOI0I
;
else
assign
CAHBLTlII0I
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTOO00
=
CAHBLTI0l0
;
else
assign
CAHBLTOO00
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTI000
=
CAHBLTlI00
;
else
assign
CAHBLTI000
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTlI10
=
CAHBLTOO10
;
else
assign
CAHBLTlI10
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTOOO1
=
CAHBLTI010
;
else
assign
CAHBLTOOO1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTI0O1
=
CAHBLTlIO1
;
else
assign
CAHBLTI0O1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTlII1
=
CAHBLTOOI1
;
else
assign
CAHBLTlII1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTOOl1
=
CAHBLTI0I1
;
else
assign
CAHBLTOOl1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTI0l1
=
CAHBLTlIl1
;
else
assign
CAHBLTI0l1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTlI01
=
CAHBLTOO01
;
else
assign
CAHBLTlI01
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTOO11
=
CAHBLTI001
;
else
assign
CAHBLTOO11
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTI011
=
CAHBLTlI11
;
else
assign
CAHBLTI011
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTlIOOI
=
CAHBLTOOOOI
;
else
assign
CAHBLTlIOOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTOOIOI
=
CAHBLTI0OOI
;
else
assign
CAHBLTOOIOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTI0IOI
=
CAHBLTlIIOI
;
else
assign
CAHBLTI0IOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTlIlOI
=
CAHBLTOOlOI
;
else
assign
CAHBLTlIlOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTOO0OI
=
CAHBLTI0lOI
;
else
assign
CAHBLTOO0OI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTI00OI
=
CAHBLTlI0OI
;
else
assign
CAHBLTI00OI
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTlI1OI
=
CAHBLTOO1OI
;
else
assign
CAHBLTlI1OI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTIOOII
=
CAHBLTl01OI
;
else
assign
CAHBLTIOOII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTl0OII
=
CAHBLTOlOII
;
else
assign
CAHBLTl0OII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTOlIII
=
CAHBLTIOIII
;
else
assign
CAHBLTOlIII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTIOlII
=
CAHBLTl0III
;
else
assign
CAHBLTIOlII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTl0lII
=
CAHBLTOllII
;
else
assign
CAHBLTl0lII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOl0II
=
CAHBLTIO0II
;
else
assign
CAHBLTOl0II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIO1II
=
CAHBLTl00II
;
else
assign
CAHBLTIO1II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTl01II
=
CAHBLTOl1II
;
else
assign
CAHBLTl01II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOlOlI
=
CAHBLTIOOlI
;
else
assign
CAHBLTOlOlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTIOIlI
=
CAHBLTl0OlI
;
else
assign
CAHBLTIOIlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTl0IlI
=
CAHBLTOlIlI
;
else
assign
CAHBLTl0IlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOlllI
=
CAHBLTIOllI
;
else
assign
CAHBLTOlllI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTIO0lI
=
CAHBLTl0llI
;
else
assign
CAHBLTIO0lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTl00lI
=
CAHBLTOl0lI
;
else
assign
CAHBLTl00lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTOl1lI
=
CAHBLTIO1lI
;
else
assign
CAHBLTOl1lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTIOO0I
=
CAHBLTl01lI
;
else
assign
CAHBLTIOO0I
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTl0O0I
=
CAHBLTOlO0I
;
else
assign
CAHBLTl0O0I
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOlI0I
=
CAHBLTIOI0I
;
else
assign
CAHBLTOlI0I
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTl0l0
=
CAHBLTOll0
;
else
assign
CAHBLTl0l0
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTOl00
=
CAHBLTIO00
;
else
assign
CAHBLTOl00
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTIO10
=
CAHBLTl000
;
else
assign
CAHBLTIO10
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTl010
=
CAHBLTOl10
;
else
assign
CAHBLTl010
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTOlO1
=
CAHBLTIOO1
;
else
assign
CAHBLTOlO1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTIOI1
=
CAHBLTl0O1
;
else
assign
CAHBLTIOI1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTl0I1
=
CAHBLTOlI1
;
else
assign
CAHBLTl0I1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTOll1
=
CAHBLTIOl1
;
else
assign
CAHBLTOll1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTIO01
=
CAHBLTl0l1
;
else
assign
CAHBLTIO01
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTl001
=
CAHBLTOl01
;
else
assign
CAHBLTl001
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTOl11
=
CAHBLTIO11
;
else
assign
CAHBLTOl11
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTIOOOI
=
CAHBLTl011
;
else
assign
CAHBLTIOOOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTl0OOI
=
CAHBLTOlOOI
;
else
assign
CAHBLTl0OOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTOlIOI
=
CAHBLTIOIOI
;
else
assign
CAHBLTOlIOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTIOlOI
=
CAHBLTl0IOI
;
else
assign
CAHBLTIOlOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTl0lOI
=
CAHBLTOllOI
;
else
assign
CAHBLTl0lOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTOl0OI
=
CAHBLTIO0OI
;
else
assign
CAHBLTOl0OI
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTIO1OI
=
CAHBLTl00OI
;
else
assign
CAHBLTIO1OI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTO11OI
=
CAHBLTIl1OI
;
else
assign
CAHBLTO11OI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTIlOII
=
CAHBLTlOOII
;
else
assign
CAHBLTIlOII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTlOIII
=
CAHBLTO1OII
;
else
assign
CAHBLTlOIII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTO1III
=
CAHBLTIlIII
;
else
assign
CAHBLTO1III
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTIllII
=
CAHBLTlOlII
;
else
assign
CAHBLTIllII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTlO0II
=
CAHBLTO1lII
;
else
assign
CAHBLTlO0II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTO10II
=
CAHBLTIl0II
;
else
assign
CAHBLTO10II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTIl1II
=
CAHBLTlO1II
;
else
assign
CAHBLTIl1II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTlOOlI
=
CAHBLTO11II
;
else
assign
CAHBLTlOOlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTO1OlI
=
CAHBLTIlOlI
;
else
assign
CAHBLTO1OlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTIlIlI
=
CAHBLTlOIlI
;
else
assign
CAHBLTIlIlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTlOllI
=
CAHBLTO1IlI
;
else
assign
CAHBLTlOllI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTO1llI
=
CAHBLTIlllI
;
else
assign
CAHBLTO1llI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTIl0lI
=
CAHBLTlO0lI
;
else
assign
CAHBLTIl0lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTlO1lI
=
CAHBLTO10lI
;
else
assign
CAHBLTlO1lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTO11lI
=
CAHBLTIl1lI
;
else
assign
CAHBLTO11lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTIlO0I
=
CAHBLTlOO0I
;
else
assign
CAHBLTIlO0I
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTlOI0I
=
CAHBLTO1O0I
;
else
assign
CAHBLTlOI0I
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTO1l0
=
CAHBLTIll0
;
else
assign
CAHBLTO1l0
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTIl00
=
CAHBLTlO00
;
else
assign
CAHBLTIl00
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTlO10
=
CAHBLTO100
;
else
assign
CAHBLTlO10
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTO110
=
CAHBLTIl10
;
else
assign
CAHBLTO110
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTIlO1
=
CAHBLTlOO1
;
else
assign
CAHBLTIlO1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTlOI1
=
CAHBLTO1O1
;
else
assign
CAHBLTlOI1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTO1I1
=
CAHBLTIlI1
;
else
assign
CAHBLTO1I1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTIll1
=
CAHBLTlOl1
;
else
assign
CAHBLTIll1
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTlO01
=
CAHBLTO1l1
;
else
assign
CAHBLTlO01
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTO101
=
CAHBLTIl01
;
else
assign
CAHBLTO101
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTIl11
=
CAHBLTlO11
;
else
assign
CAHBLTIl11
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTlOOOI
=
CAHBLTO111
;
else
assign
CAHBLTlOOOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTO1OOI
=
CAHBLTIlOOI
;
else
assign
CAHBLTO1OOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTIlIOI
=
CAHBLTlOIOI
;
else
assign
CAHBLTIlIOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTlOlOI
=
CAHBLTO1IOI
;
else
assign
CAHBLTlOlOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTO1lOI
=
CAHBLTIllOI
;
else
assign
CAHBLTO1lOI
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTIl0OI
=
CAHBLTlO0OI
;
else
assign
CAHBLTIl0OI
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTlO1OI
=
CAHBLTO10OI
;
else
assign
CAHBLTlO1OI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTI11OI
=
CAHBLTll1OI
;
else
assign
CAHBLTI11OI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTllOII
=
CAHBLTOIOII
;
else
assign
CAHBLTllOII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTOIIII
=
CAHBLTI1OII
;
else
assign
CAHBLTOIIII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTI1III
=
CAHBLTllIII
;
else
assign
CAHBLTI1III
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTlllII
=
CAHBLTOIlII
;
else
assign
CAHBLTlllII
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOI0II
=
CAHBLTI1lII
;
else
assign
CAHBLTOI0II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTI10II
=
CAHBLTll0II
;
else
assign
CAHBLTI10II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTll1II
=
CAHBLTOI1II
;
else
assign
CAHBLTll1II
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOIOlI
=
CAHBLTI11II
;
else
assign
CAHBLTOIOlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTI1OlI
=
CAHBLTllOlI
;
else
assign
CAHBLTI1OlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTllIlI
=
CAHBLTOIIlI
;
else
assign
CAHBLTllIlI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOIllI
=
CAHBLTI1IlI
;
else
assign
CAHBLTOIllI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTI1llI
=
CAHBLTllllI
;
else
assign
CAHBLTI1llI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTll0lI
=
CAHBLTOI0lI
;
else
assign
CAHBLTll0lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTOI1lI
=
CAHBLTI10lI
;
else
assign
CAHBLTOI1lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTI11lI
=
CAHBLTll1lI
;
else
assign
CAHBLTI11lI
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTllO0I
=
CAHBLTOIO0I
;
else
assign
CAHBLTllO0I
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOII0I
=
CAHBLTI1O0I
;
else
assign
CAHBLTOII0I
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTI1OOl
=
CAHBLTOlll
;
else
assign
CAHBLTI1OOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTl1OOl
=
CAHBLTOlll
;
else
assign
CAHBLTl1OOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTOOIOl
=
CAHBLTOlll
;
else
assign
CAHBLTOOIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTIOIOl
=
CAHBLTOlll
;
else
assign
CAHBLTIOIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTlOIOl
=
CAHBLTOlll
;
else
assign
CAHBLTlOIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTOIIOl
=
CAHBLTOlll
;
else
assign
CAHBLTOIIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTIIIOl
=
CAHBLTOlll
;
else
assign
CAHBLTIIIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTlIIOl
=
CAHBLTOlll
;
else
assign
CAHBLTlIIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTOlIOl
=
CAHBLTOlll
;
else
assign
CAHBLTOlIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTIlIOl
=
CAHBLTOlll
;
else
assign
CAHBLTIlIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTllIOl
=
CAHBLTOlll
;
else
assign
CAHBLTllIOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTO0IOl
=
CAHBLTOlll
;
else
assign
CAHBLTO0IOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTI0IOl
=
CAHBLTOlll
;
else
assign
CAHBLTI0IOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTl0IOl
=
CAHBLTOlll
;
else
assign
CAHBLTl0IOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTO1IOl
=
CAHBLTOlll
;
else
assign
CAHBLTO1IOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTI1IOl
=
CAHBLTOlll
;
else
assign
CAHBLTI1IOl
=
32
'h
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTl1IOl
=
CAHBLTOlll
;
else
assign
CAHBLTl1IOl
=
32
'h
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOOlOl
=
CAHBLTOlll
;
else
assign
CAHBLTOOlOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTIOlOl
=
CAHBLTI0ll
;
else
assign
CAHBLTIOlOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTlOlOl
=
CAHBLTI0ll
;
else
assign
CAHBLTlOlOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTOIlOl
=
CAHBLTI0ll
;
else
assign
CAHBLTOIlOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTIIlOl
=
CAHBLTI0ll
;
else
assign
CAHBLTIIlOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTlIlOl
=
CAHBLTI0ll
;
else
assign
CAHBLTlIlOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOllOl
=
CAHBLTI0ll
;
else
assign
CAHBLTOllOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIllOl
=
CAHBLTI0ll
;
else
assign
CAHBLTIllOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTlllOl
=
CAHBLTI0ll
;
else
assign
CAHBLTlllOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTO0lOl
=
CAHBLTI0ll
;
else
assign
CAHBLTO0lOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTI0lOl
=
CAHBLTI0ll
;
else
assign
CAHBLTI0lOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTl0lOl
=
CAHBLTI0ll
;
else
assign
CAHBLTl0lOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTO1lOl
=
CAHBLTI0ll
;
else
assign
CAHBLTO1lOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTI1lOl
=
CAHBLTI0ll
;
else
assign
CAHBLTI1lOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTl1lOl
=
CAHBLTI0ll
;
else
assign
CAHBLTl1lOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTOO0Ol
=
CAHBLTI0ll
;
else
assign
CAHBLTOO0Ol
=
32
'h
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTIO0Ol
=
CAHBLTI0ll
;
else
assign
CAHBLTIO0Ol
=
32
'h
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTlO0Ol
=
CAHBLTI0ll
;
else
assign
CAHBLTlO0Ol
=
32
'h
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOI0Ol
=
CAHBLTI0ll
;
else
assign
CAHBLTOI0Ol
=
32
'h
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTI0OIl
=
CAHBLTll1
;
else
assign
CAHBLTI0OIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTl0OIl
=
CAHBLTll1
;
else
assign
CAHBLTl0OIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTO1OIl
=
CAHBLTll1
;
else
assign
CAHBLTO1OIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTI1OIl
=
CAHBLTll1
;
else
assign
CAHBLTI1OIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTl1OIl
=
CAHBLTll1
;
else
assign
CAHBLTl1OIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTOOIIl
=
CAHBLTll1
;
else
assign
CAHBLTOOIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTIOIIl
=
CAHBLTll1
;
else
assign
CAHBLTIOIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTlOIIl
=
CAHBLTll1
;
else
assign
CAHBLTlOIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTOIIIl
=
CAHBLTll1
;
else
assign
CAHBLTOIIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTIIIIl
=
CAHBLTll1
;
else
assign
CAHBLTIIIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTlIIIl
=
CAHBLTll1
;
else
assign
CAHBLTlIIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTOlIIl
=
CAHBLTll1
;
else
assign
CAHBLTOlIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTIlIIl
=
CAHBLTll1
;
else
assign
CAHBLTIlIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTllIIl
=
CAHBLTll1
;
else
assign
CAHBLTllIIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTO0IIl
=
CAHBLTll1
;
else
assign
CAHBLTO0IIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTI0IIl
=
CAHBLTll1
;
else
assign
CAHBLTI0IIl
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTl0IIl
=
CAHBLTll1
;
else
assign
CAHBLTl0IIl
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTO1IIl
=
CAHBLTll1
;
else
assign
CAHBLTO1IIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTI1IIl
=
CAHBLTO01
;
else
assign
CAHBLTI1IIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTl1IIl
=
CAHBLTO01
;
else
assign
CAHBLTl1IIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTOOlIl
=
CAHBLTO01
;
else
assign
CAHBLTOOlIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTIOlIl
=
CAHBLTO01
;
else
assign
CAHBLTIOlIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTlOlIl
=
CAHBLTO01
;
else
assign
CAHBLTlOlIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOIlIl
=
CAHBLTO01
;
else
assign
CAHBLTOIlIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIIlIl
=
CAHBLTO01
;
else
assign
CAHBLTIIlIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTlIlIl
=
CAHBLTO01
;
else
assign
CAHBLTlIlIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOllIl
=
CAHBLTO01
;
else
assign
CAHBLTOllIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTIllIl
=
CAHBLTO01
;
else
assign
CAHBLTIllIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTlllIl
=
CAHBLTO01
;
else
assign
CAHBLTlllIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTO0lIl
=
CAHBLTO01
;
else
assign
CAHBLTO0lIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTI0lIl
=
CAHBLTO01
;
else
assign
CAHBLTI0lIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTl0lIl
=
CAHBLTO01
;
else
assign
CAHBLTl0lIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTO1lIl
=
CAHBLTO01
;
else
assign
CAHBLTO1lIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTI1lIl
=
CAHBLTO01
;
else
assign
CAHBLTI1lIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTl1lIl
=
CAHBLTO01
;
else
assign
CAHBLTl1lIl
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOO0Il
=
CAHBLTO01
;
else
assign
CAHBLTOO0Il
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTII0Ol
=
CAHBLTIlll
;
else
assign
CAHBLTII0Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTlI0Ol
=
CAHBLTIlll
;
else
assign
CAHBLTlI0Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTOl0Ol
=
CAHBLTIlll
;
else
assign
CAHBLTOl0Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTIl0Ol
=
CAHBLTIlll
;
else
assign
CAHBLTIl0Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTll0Ol
=
CAHBLTIlll
;
else
assign
CAHBLTll0Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTO00Ol
=
CAHBLTIlll
;
else
assign
CAHBLTO00Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTI00Ol
=
CAHBLTIlll
;
else
assign
CAHBLTI00Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTl00Ol
=
CAHBLTIlll
;
else
assign
CAHBLTl00Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTO10Ol
=
CAHBLTIlll
;
else
assign
CAHBLTO10Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTI10Ol
=
CAHBLTIlll
;
else
assign
CAHBLTI10Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTl10Ol
=
CAHBLTIlll
;
else
assign
CAHBLTl10Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTOO1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTOO1Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTIO1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTIO1Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTlO1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTlO1Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTOI1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTOI1Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTII1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTII1Ol
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTlI1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTlI1Ol
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOl1Ol
=
CAHBLTIlll
;
else
assign
CAHBLTOl1Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTIl1Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTIl1Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTll1Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTll1Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTO01Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTO01Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTI01Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTI01Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTl01Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTl01Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTO11Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTO11Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTI11Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTI11Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTl11Ol
=
CAHBLTl0ll
;
else
assign
CAHBLTl11Ol
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOOOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTOOOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTIOOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTIOOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTlOOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTlOOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOIOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTOIOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTIIOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTIIOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTlIOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTlIOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTOlOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTOlOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTIlOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTIlOIl
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTllOIl
=
CAHBLTl0ll
;
else
assign
CAHBLTllOIl
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTO0OIl
=
CAHBLTl0ll
;
else
assign
CAHBLTO0OIl
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTIO0Il
=
CAHBLTllll
;
else
assign
CAHBLTIO0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTlO0Il
=
CAHBLTllll
;
else
assign
CAHBLTlO0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTOI0Il
=
CAHBLTllll
;
else
assign
CAHBLTOI0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTII0Il
=
CAHBLTllll
;
else
assign
CAHBLTII0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTlI0Il
=
CAHBLTllll
;
else
assign
CAHBLTlI0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTOl0Il
=
CAHBLTllll
;
else
assign
CAHBLTOl0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTIl0Il
=
CAHBLTllll
;
else
assign
CAHBLTIl0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTll0Il
=
CAHBLTllll
;
else
assign
CAHBLTll0Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTO00Il
=
CAHBLTllll
;
else
assign
CAHBLTO00Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTI00Il
=
CAHBLTllll
;
else
assign
CAHBLTI00Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTl00Il
=
CAHBLTllll
;
else
assign
CAHBLTl00Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTO10Il
=
CAHBLTllll
;
else
assign
CAHBLTO10Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTI10Il
=
CAHBLTllll
;
else
assign
CAHBLTI10Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTl10Il
=
CAHBLTllll
;
else
assign
CAHBLTl10Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTOO1Il
=
CAHBLTllll
;
else
assign
CAHBLTOO1Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTIO1Il
=
CAHBLTllll
;
else
assign
CAHBLTIO1Il
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTlO1Il
=
CAHBLTllll
;
else
assign
CAHBLTlO1Il
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOI1Il
=
CAHBLTllll
;
else
assign
CAHBLTOI1Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTII1Il
=
CAHBLTO1ll
;
else
assign
CAHBLTII1Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTlI1Il
=
CAHBLTO1ll
;
else
assign
CAHBLTlI1Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTOl1Il
=
CAHBLTO1ll
;
else
assign
CAHBLTOl1Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTIl1Il
=
CAHBLTO1ll
;
else
assign
CAHBLTIl1Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTll1Il
=
CAHBLTO1ll
;
else
assign
CAHBLTll1Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTO01Il
=
CAHBLTO1ll
;
else
assign
CAHBLTO01Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTI01Il
=
CAHBLTO1ll
;
else
assign
CAHBLTI01Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTl01Il
=
CAHBLTO1ll
;
else
assign
CAHBLTl01Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTO11Il
=
CAHBLTO1ll
;
else
assign
CAHBLTO11Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTI11Il
=
CAHBLTO1ll
;
else
assign
CAHBLTI11Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTl11Il
=
CAHBLTO1ll
;
else
assign
CAHBLTl11Il
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOOOll
=
CAHBLTO1ll
;
else
assign
CAHBLTOOOll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTIOOll
=
CAHBLTO1ll
;
else
assign
CAHBLTIOOll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTlOOll
=
CAHBLTO1ll
;
else
assign
CAHBLTlOOll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTOIOll
=
CAHBLTO1ll
;
else
assign
CAHBLTOIOll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTIIOll
=
CAHBLTO1ll
;
else
assign
CAHBLTIIOll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTlIOll
=
CAHBLTO1ll
;
else
assign
CAHBLTlIOll
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOlOll
=
CAHBLTO1ll
;
else
assign
CAHBLTOlOll
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTIlOll
=
CAHBLTO0ll
;
else
assign
CAHBLTIlOll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTllOll
=
CAHBLTO0ll
;
else
assign
CAHBLTllOll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTO0Oll
=
CAHBLTO0ll
;
else
assign
CAHBLTO0Oll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTI0Oll
=
CAHBLTO0ll
;
else
assign
CAHBLTI0Oll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTl0Oll
=
CAHBLTO0ll
;
else
assign
CAHBLTl0Oll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTO1Oll
=
CAHBLTO0ll
;
else
assign
CAHBLTO1Oll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTI1Oll
=
CAHBLTO0ll
;
else
assign
CAHBLTI1Oll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTl1Oll
=
CAHBLTO0ll
;
else
assign
CAHBLTl1Oll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTOOIll
=
CAHBLTO0ll
;
else
assign
CAHBLTOOIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTIOIll
=
CAHBLTO0ll
;
else
assign
CAHBLTIOIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTlOIll
=
CAHBLTO0ll
;
else
assign
CAHBLTlOIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTOIIll
=
CAHBLTO0ll
;
else
assign
CAHBLTOIIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTIIIll
=
CAHBLTO0ll
;
else
assign
CAHBLTIIIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTlIIll
=
CAHBLTO0ll
;
else
assign
CAHBLTlIIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTOlIll
=
CAHBLTO0ll
;
else
assign
CAHBLTOlIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTIlIll
=
CAHBLTO0ll
;
else
assign
CAHBLTIlIll
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTllIll
=
CAHBLTO0ll
;
else
assign
CAHBLTllIll
=
1
'b
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTO0Ill
=
CAHBLTO0ll
;
else
assign
CAHBLTO0Ill
=
1
'b
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTI0Ill
=
CAHBLTI1ll
;
else
assign
CAHBLTI0Ill
=
1
'b
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTl0Ill
=
CAHBLTI1ll
;
else
assign
CAHBLTl0Ill
=
1
'b
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTO1Ill
=
CAHBLTI1ll
;
else
assign
CAHBLTO1Ill
=
1
'b
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTI1Ill
=
CAHBLTI1ll
;
else
assign
CAHBLTI1Ill
=
1
'b
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTl1Ill
=
CAHBLTI1ll
;
else
assign
CAHBLTl1Ill
=
1
'b
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOOlll
=
CAHBLTI1ll
;
else
assign
CAHBLTOOlll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIOlll
=
CAHBLTI1ll
;
else
assign
CAHBLTIOlll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTlOlll
=
CAHBLTI1ll
;
else
assign
CAHBLTlOlll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOIlll
=
CAHBLTI1ll
;
else
assign
CAHBLTOIlll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTIIlll
=
CAHBLTI1ll
;
else
assign
CAHBLTIIlll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTlIlll
=
CAHBLTI1ll
;
else
assign
CAHBLTlIlll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOllll
=
CAHBLTI1ll
;
else
assign
CAHBLTOllll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTIllll
=
CAHBLTI1ll
;
else
assign
CAHBLTIllll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTlllll
=
CAHBLTI1ll
;
else
assign
CAHBLTlllll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTO0lll
=
CAHBLTI1ll
;
else
assign
CAHBLTO0lll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTI0lll
=
CAHBLTI1ll
;
else
assign
CAHBLTI0lll
=
1
'b
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTl0lll
=
CAHBLTI1ll
;
else
assign
CAHBLTl0lll
=
1
'b
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTO1lll
=
CAHBLTI1ll
;
else
assign
CAHBLTO1lll
=
1
'b
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTI1lll
=
CAHBLTlIl0
;
else
assign
CAHBLTI1lll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTl1lll
=
CAHBLTlIl0
;
else
assign
CAHBLTl1lll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTOO0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTOO0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTIO0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTIO0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTlO0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTlO0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTOI0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTOI0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTII0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTII0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTlI0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTlI0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTOl0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTOl0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTIl0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTIl0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTll0ll
=
CAHBLTlIl0
;
else
assign
CAHBLTll0ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTO00ll
=
CAHBLTlIl0
;
else
assign
CAHBLTO00ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTI00ll
=
CAHBLTlIl0
;
else
assign
CAHBLTI00ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTl00ll
=
CAHBLTlIl0
;
else
assign
CAHBLTl00ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTO10ll
=
CAHBLTlIl0
;
else
assign
CAHBLTO10ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTI10ll
=
CAHBLTlIl0
;
else
assign
CAHBLTI10ll
=
1
'b
1
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTl10ll
=
CAHBLTlIl0
;
else
assign
CAHBLTl10ll
=
1
'b
1
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOO1ll
=
CAHBLTlIl0
;
else
assign
CAHBLTOO1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTIO1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTIO1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTlO1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTlO1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTOI1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTOI1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTII1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTII1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTlI1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTlI1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOl1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTOl1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIl1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTIl1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTll1ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTll1ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTO01ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTO01ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTI01ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTI01ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTl01ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTl01ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTO11ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTO11ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTI11ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTI11ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTl11ll
=
CAHBLTOl1OI
;
else
assign
CAHBLTl11ll
=
1
'b
1
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTOOO0l
=
CAHBLTOl1OI
;
else
assign
CAHBLTOOO0l
=
1
'b
1
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTIOO0l
=
CAHBLTOl1OI
;
else
assign
CAHBLTIOO0l
=
1
'b
1
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTlOO0l
=
CAHBLTOl1OI
;
else
assign
CAHBLTlOO0l
=
1
'b
1
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTOIO0l
=
CAHBLTOl1OI
;
else
assign
CAHBLTOIO0l
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTllI0I
=
HRDATA_S0
;
else
assign
CAHBLTllI0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTO0I0I
=
HRDATA_S1
;
else
assign
CAHBLTO0I0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTI0I0I
=
HRDATA_S2
;
else
assign
CAHBLTI0I0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTl0I0I
=
HRDATA_S3
;
else
assign
CAHBLTl0I0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTO1I0I
=
HRDATA_S4
;
else
assign
CAHBLTO1I0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTI1I0I
=
HRDATA_S5
;
else
assign
CAHBLTI1I0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTl1I0I
=
HRDATA_S6
;
else
assign
CAHBLTl1I0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTOOl0I
=
HRDATA_S7
;
else
assign
CAHBLTOOl0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTIOl0I
=
HRDATA_S8
;
else
assign
CAHBLTIOl0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTlOl0I
=
HRDATA_S9
;
else
assign
CAHBLTlOl0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTOIl0I
=
HRDATA_S10
;
else
assign
CAHBLTOIl0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTIIl0I
=
HRDATA_S11
;
else
assign
CAHBLTIIl0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTlIl0I
=
HRDATA_S12
;
else
assign
CAHBLTlIl0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTOll0I
=
HRDATA_S13
;
else
assign
CAHBLTOll0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTIll0I
=
HRDATA_S14
;
else
assign
CAHBLTIll0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTlll0I
=
HRDATA_S15
;
else
assign
CAHBLTlll0I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTO0l0I
=
HRDATA_SHG
;
else
assign
CAHBLTO0l0I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTI0l0I
=
HRDATA_S0
;
else
assign
CAHBLTI0l0I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTl0l0I
=
HRDATA_S1
;
else
assign
CAHBLTl0l0I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTO1l0I
=
HRDATA_S2
;
else
assign
CAHBLTO1l0I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTI1l0I
=
HRDATA_S3
;
else
assign
CAHBLTI1l0I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTl1l0I
=
HRDATA_S4
;
else
assign
CAHBLTl1l0I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOO00I
=
HRDATA_S5
;
else
assign
CAHBLTOO00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIO00I
=
HRDATA_S6
;
else
assign
CAHBLTIO00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTlO00I
=
HRDATA_S7
;
else
assign
CAHBLTlO00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOI00I
=
HRDATA_S8
;
else
assign
CAHBLTOI00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTII00I
=
HRDATA_S9
;
else
assign
CAHBLTII00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTlI00I
=
HRDATA_S10
;
else
assign
CAHBLTlI00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOl00I
=
HRDATA_S11
;
else
assign
CAHBLTOl00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTIl00I
=
HRDATA_S12
;
else
assign
CAHBLTIl00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTll00I
=
HRDATA_S13
;
else
assign
CAHBLTll00I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTO000I
=
HRDATA_S14
;
else
assign
CAHBLTO000I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTI000I
=
HRDATA_S15
;
else
assign
CAHBLTI000I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTl000I
=
HRDATA_SHG
;
else
assign
CAHBLTl000I
=
32
'h
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTIl01I
=
HWDATA_M0
;
else
assign
CAHBLTIl01I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTll01I
=
HWDATA_M0
;
else
assign
CAHBLTll01I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTO001I
=
HWDATA_M0
;
else
assign
CAHBLTO001I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTI001I
=
HWDATA_M0
;
else
assign
CAHBLTI001I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTl001I
=
HWDATA_M0
;
else
assign
CAHBLTl001I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTO101I
=
HWDATA_M0
;
else
assign
CAHBLTO101I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTI101I
=
HWDATA_M0
;
else
assign
CAHBLTI101I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTl101I
=
HWDATA_M0
;
else
assign
CAHBLTl101I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTOO11I
=
HWDATA_M0
;
else
assign
CAHBLTOO11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTIO11I
=
HWDATA_M0
;
else
assign
CAHBLTIO11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTlO11I
=
HWDATA_M0
;
else
assign
CAHBLTlO11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTOI11I
=
HWDATA_M0
;
else
assign
CAHBLTOI11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTII11I
=
HWDATA_M0
;
else
assign
CAHBLTII11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTlI11I
=
HWDATA_M0
;
else
assign
CAHBLTlI11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTOl11I
=
HWDATA_M0
;
else
assign
CAHBLTOl11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTIl11I
=
HWDATA_M0
;
else
assign
CAHBLTIl11I
=
32
'h
0
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTll11I
=
HWDATA_M0
;
else
assign
CAHBLTll11I
=
32
'h
0
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTO011I
=
HWDATA_M0
;
else
assign
CAHBLTO011I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTI011I
=
HWDATA_M1
;
else
assign
CAHBLTI011I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTl011I
=
HWDATA_M1
;
else
assign
CAHBLTl011I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTO111I
=
HWDATA_M1
;
else
assign
CAHBLTO111I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTI111I
=
HWDATA_M1
;
else
assign
CAHBLTI111I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTl111I
=
HWDATA_M1
;
else
assign
CAHBLTl111I
=
32
'h
0
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTOOOOl
=
HWDATA_M1
;
else
assign
CAHBLTOOOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTIOOOl
=
HWDATA_M1
;
else
assign
CAHBLTIOOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTlOOOl
=
HWDATA_M1
;
else
assign
CAHBLTlOOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTOIOOl
=
HWDATA_M1
;
else
assign
CAHBLTOIOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTIIOOl
=
HWDATA_M1
;
else
assign
CAHBLTIIOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTlIOOl
=
HWDATA_M1
;
else
assign
CAHBLTlIOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTOlOOl
=
HWDATA_M1
;
else
assign
CAHBLTOlOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTIlOOl
=
HWDATA_M1
;
else
assign
CAHBLTIlOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTllOOl
=
HWDATA_M1
;
else
assign
CAHBLTllOOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTO0OOl
=
HWDATA_M1
;
else
assign
CAHBLTO0OOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTI0OOl
=
HWDATA_M1
;
else
assign
CAHBLTI0OOl
=
32
'h
0
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTl0OOl
=
HWDATA_M1
;
else
assign
CAHBLTl0OOl
=
32
'h
0
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTO1OOl
=
HWDATA_M1
;
else
assign
CAHBLTO1OOl
=
32
'h
0
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
)
assign
CAHBLTO100I
=
HREADYOUT_S0
;
else
assign
CAHBLTO100I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
1
]
)
assign
CAHBLTI100I
=
HREADYOUT_S1
;
else
assign
CAHBLTI100I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
2
]
)
assign
CAHBLTl100I
=
HREADYOUT_S2
;
else
assign
CAHBLTl100I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
3
]
)
assign
CAHBLTOO10I
=
HREADYOUT_S3
;
else
assign
CAHBLTOO10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
4
]
)
assign
CAHBLTIO10I
=
HREADYOUT_S4
;
else
assign
CAHBLTIO10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
5
]
)
assign
CAHBLTlO10I
=
HREADYOUT_S5
;
else
assign
CAHBLTlO10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
6
]
)
assign
CAHBLTOI10I
=
HREADYOUT_S6
;
else
assign
CAHBLTOI10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
7
]
)
assign
CAHBLTII10I
=
HREADYOUT_S7
;
else
assign
CAHBLTII10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
8
]
)
assign
CAHBLTlI10I
=
HREADYOUT_S8
;
else
assign
CAHBLTlI10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
9
]
)
assign
CAHBLTOl10I
=
HREADYOUT_S9
;
else
assign
CAHBLTOl10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
10
]
)
assign
CAHBLTIl10I
=
HREADYOUT_S10
;
else
assign
CAHBLTIl10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
11
]
)
assign
CAHBLTll10I
=
HREADYOUT_S11
;
else
assign
CAHBLTll10I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
12
]
)
assign
CAHBLTO010I
=
HREADYOUT_S12
;
else
assign
CAHBLTO010I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
13
]
)
assign
CAHBLTI010I
=
HREADYOUT_S13
;
else
assign
CAHBLTI010I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
14
]
)
assign
CAHBLTl010I
=
HREADYOUT_S14
;
else
assign
CAHBLTl010I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
15
]
)
assign
CAHBLTO110I
=
HREADYOUT_S15
;
else
assign
CAHBLTO110I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
16
]
)
assign
CAHBLTI110I
=
HREADYOUT_SHG
;
else
assign
CAHBLTI110I
=
1
'b
1
;
if
(
CAHBLTO0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTl110I
=
CAHBLTIlI0I
;
else
assign
CAHBLTl110I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
0
]
)
assign
CAHBLTOOO1I
=
HREADYOUT_S0
;
else
assign
CAHBLTOOO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
1
]
)
assign
CAHBLTIOO1I
=
HREADYOUT_S1
;
else
assign
CAHBLTIOO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
2
]
)
assign
CAHBLTlOO1I
=
HREADYOUT_S2
;
else
assign
CAHBLTlOO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
3
]
)
assign
CAHBLTOIO1I
=
HREADYOUT_S3
;
else
assign
CAHBLTOIO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
4
]
)
assign
CAHBLTIIO1I
=
HREADYOUT_S4
;
else
assign
CAHBLTIIO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
5
]
)
assign
CAHBLTlIO1I
=
HREADYOUT_S5
;
else
assign
CAHBLTlIO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
6
]
)
assign
CAHBLTOlO1I
=
HREADYOUT_S6
;
else
assign
CAHBLTOlO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
7
]
)
assign
CAHBLTIlO1I
=
HREADYOUT_S7
;
else
assign
CAHBLTIlO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
8
]
)
assign
CAHBLTllO1I
=
HREADYOUT_S8
;
else
assign
CAHBLTllO1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
9
]
)
assign
CAHBLTO0O1I
=
HREADYOUT_S9
;
else
assign
CAHBLTO0O1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
10
]
)
assign
CAHBLTI0O1I
=
HREADYOUT_S10
;
else
assign
CAHBLTI0O1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
11
]
)
assign
CAHBLTl0O1I
=
HREADYOUT_S11
;
else
assign
CAHBLTl0O1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
12
]
)
assign
CAHBLTO1O1I
=
HREADYOUT_S12
;
else
assign
CAHBLTO1O1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
13
]
)
assign
CAHBLTI1O1I
=
HREADYOUT_S13
;
else
assign
CAHBLTI1O1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
14
]
)
assign
CAHBLTl1O1I
=
HREADYOUT_S14
;
else
assign
CAHBLTl1O1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
15
]
)
assign
CAHBLTOOI1I
=
HREADYOUT_S15
;
else
assign
CAHBLTOOI1I
=
1
'b
1
;
if
(
CAHBLTIIl0
[
16
]
)
assign
CAHBLTIOI1I
=
HREADYOUT_SHG
;
else
assign
CAHBLTIOI1I
=
1
'b
1
;
if
(
CAHBLTI0O0
[
15
:
0
]
!=
0
)
assign
CAHBLTlOI1I
=
CAHBLTIlI0I
;
else
assign
CAHBLTlOI1I
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
|
CAHBLTIIl0
[
0
]
)
assign
CAHBLTOII1I
=
HREADYOUT_S0
;
else
assign
CAHBLTOII1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
1
]
|
CAHBLTIIl0
[
1
]
)
assign
CAHBLTIII1I
=
HREADYOUT_S1
;
else
assign
CAHBLTIII1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
2
]
|
CAHBLTIIl0
[
2
]
)
assign
CAHBLTlII1I
=
HREADYOUT_S2
;
else
assign
CAHBLTlII1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
3
]
|
CAHBLTIIl0
[
3
]
)
assign
CAHBLTOlI1I
=
HREADYOUT_S3
;
else
assign
CAHBLTOlI1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
4
]
|
CAHBLTIIl0
[
4
]
)
assign
CAHBLTIlI1I
=
HREADYOUT_S4
;
else
assign
CAHBLTIlI1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
5
]
|
CAHBLTIIl0
[
5
]
)
assign
CAHBLTllI1I
=
HREADYOUT_S5
;
else
assign
CAHBLTllI1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
6
]
|
CAHBLTIIl0
[
6
]
)
assign
CAHBLTO0I1I
=
HREADYOUT_S6
;
else
assign
CAHBLTO0I1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
7
]
|
CAHBLTIIl0
[
7
]
)
assign
CAHBLTI0I1I
=
HREADYOUT_S7
;
else
assign
CAHBLTI0I1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
8
]
|
CAHBLTIIl0
[
8
]
)
assign
CAHBLTl0I1I
=
HREADYOUT_S8
;
else
assign
CAHBLTl0I1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
9
]
|
CAHBLTIIl0
[
9
]
)
assign
CAHBLTO1I1I
=
HREADYOUT_S9
;
else
assign
CAHBLTO1I1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
10
]
|
CAHBLTIIl0
[
10
]
)
assign
CAHBLTI1I1I
=
HREADYOUT_S10
;
else
assign
CAHBLTI1I1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
11
]
|
CAHBLTIIl0
[
11
]
)
assign
CAHBLTl1I1I
=
HREADYOUT_S11
;
else
assign
CAHBLTl1I1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
12
]
|
CAHBLTIIl0
[
12
]
)
assign
CAHBLTOOl1I
=
HREADYOUT_S12
;
else
assign
CAHBLTOOl1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
13
]
|
CAHBLTIIl0
[
13
]
)
assign
CAHBLTIOl1I
=
HREADYOUT_S13
;
else
assign
CAHBLTIOl1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
14
]
|
CAHBLTIIl0
[
14
]
)
assign
CAHBLTlOl1I
=
HREADYOUT_S14
;
else
assign
CAHBLTlOl1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
15
]
|
CAHBLTIIl0
[
15
]
)
assign
CAHBLTOIl1I
=
HREADYOUT_S15
;
else
assign
CAHBLTOIl1I
=
1
'b
1
;
if
(
CAHBLTOIl0
[
16
]
|
CAHBLTIIl0
[
16
]
)
assign
CAHBLTIIl1I
=
HREADYOUT_SHG
;
else
assign
CAHBLTIIl1I
=
1
'b
1
;
endgenerate
generate
if
(
CAHBLTOIl0
[
0
]
|
CAHBLTIIl0
[
0
]
)
assign
CAHBLTlIl1I
=
HRESP_S0
;
else
assign
CAHBLTlIl1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
1
]
|
CAHBLTIIl0
[
1
]
)
assign
CAHBLTOll1I
=
HRESP_S1
;
else
assign
CAHBLTOll1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
2
]
|
CAHBLTIIl0
[
2
]
)
assign
CAHBLTIll1I
=
HRESP_S2
;
else
assign
CAHBLTIll1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
3
]
|
CAHBLTIIl0
[
3
]
)
assign
CAHBLTlll1I
=
HRESP_S3
;
else
assign
CAHBLTlll1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
4
]
|
CAHBLTIIl0
[
4
]
)
assign
CAHBLTO0l1I
=
HRESP_S4
;
else
assign
CAHBLTO0l1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
5
]
|
CAHBLTIIl0
[
5
]
)
assign
CAHBLTI0l1I
=
HRESP_S5
;
else
assign
CAHBLTI0l1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
6
]
|
CAHBLTIIl0
[
6
]
)
assign
CAHBLTl0l1I
=
HRESP_S6
;
else
assign
CAHBLTl0l1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
7
]
|
CAHBLTIIl0
[
7
]
)
assign
CAHBLTO1l1I
=
HRESP_S7
;
else
assign
CAHBLTO1l1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
8
]
|
CAHBLTIIl0
[
8
]
)
assign
CAHBLTI1l1I
=
HRESP_S8
;
else
assign
CAHBLTI1l1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
9
]
|
CAHBLTIIl0
[
9
]
)
assign
CAHBLTl1l1I
=
HRESP_S9
;
else
assign
CAHBLTl1l1I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
10
]
|
CAHBLTIIl0
[
10
]
)
assign
CAHBLTOO01I
=
HRESP_S10
;
else
assign
CAHBLTOO01I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
11
]
|
CAHBLTIIl0
[
11
]
)
assign
CAHBLTIO01I
=
HRESP_S11
;
else
assign
CAHBLTIO01I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
12
]
|
CAHBLTIIl0
[
12
]
)
assign
CAHBLTlO01I
=
HRESP_S12
;
else
assign
CAHBLTlO01I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
13
]
|
CAHBLTIIl0
[
13
]
)
assign
CAHBLTOI01I
=
HRESP_S13
;
else
assign
CAHBLTOI01I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
14
]
|
CAHBLTIIl0
[
14
]
)
assign
CAHBLTII01I
=
HRESP_S14
;
else
assign
CAHBLTII01I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
15
]
|
CAHBLTIIl0
[
15
]
)
assign
CAHBLTlI01I
=
HRESP_S15
;
else
assign
CAHBLTlI01I
=
1
'b
0
;
if
(
CAHBLTOIl0
[
16
]
|
CAHBLTIIl0
[
16
]
)
assign
CAHBLTOl01I
=
HRESP_SHG
;
else
assign
CAHBLTOl01I
=
1
'b
0
;
endgenerate
CAHBLTO0OI
#
(
.MODE_CFG
(
MODE_CFG
)
,
.CAHBLTI
(
CAHBLTOIl0
)
,
.CAHBLTl
(
CAHBLTO0O0
)
)
CAHBLTOlO0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTI0OI
(
HADDR_M0
)
,
.CAHBLTl0OI
(
HMASTLOCK_M0
)
,
.CAHBLTO1OI
(
HSIZE_M0
)
,
.CAHBLTI1OI
(
HTRANS_M0
)
,
.CAHBLTl1OI
(
HWRITE_M0
)
,
.CAHBLTII
(
REMAP_M0
)
,
.CAHBLTOOII
(
HRESP_M0
)
,
.CAHBLTIOII
(
HRDATA_M0
)
,
.CAHBLTlOII
(
CAHBLTIIO0l
)
,
.CAHBLTOIII
(
{
CAHBLTll0OI
,
CAHBLTI1lOI
,
CAHBLTOIlOI
,
CAHBLTllIOI
,
CAHBLTI1OOI
,
CAHBLTOIOOI
,
CAHBLTll11
,
CAHBLTI101
,
CAHBLTOI01
,
CAHBLTlll1
,
CAHBLTI1I1
,
CAHBLTOII1
,
CAHBLTllO1
,
CAHBLTI110
,
CAHBLTOI10
,
CAHBLTll00
,
CAHBLTI1l0
}
)
,
.CAHBLTIIII
(
{
CAHBLTO00OI
,
CAHBLTl1lOI
,
CAHBLTIIlOI
,
CAHBLTO0IOI
,
CAHBLTl1OOI
,
CAHBLTIIOOI
,
CAHBLTO011
,
CAHBLTl101
,
CAHBLTII01
,
CAHBLTO0l1
,
CAHBLTl1I1
,
CAHBLTIII1
,
CAHBLTO0O1
,
CAHBLTl110
,
CAHBLTII10
,
CAHBLTO000
,
CAHBLTl1l0
}
)
,
.CAHBLTlIII
(
{
CAHBLTI00OI
,
CAHBLTOO0OI
,
CAHBLTlIlOI
,
CAHBLTI0IOI
,
CAHBLTOOIOI
,
CAHBLTlIOOI
,
CAHBLTI011
,
CAHBLTOO11
,
CAHBLTlI01
,
CAHBLTI0l1
,
CAHBLTOOl1
,
CAHBLTlII1
,
CAHBLTI0O1
,
CAHBLTOOO1
,
CAHBLTlI10
,
CAHBLTI000
,
CAHBLTOO00
}
)
,
.CAHBLTOlII
(
CAHBLTOI1OI
)
,
.CAHBLTIlII
(
CAHBLTII1OI
)
,
.CAHBLTllII
(
CAHBLTlI1OI
)
,
.CAHBLTO0II
(
CAHBLTOlll
)
,
.CAHBLTI0II
(
CAHBLTll1
)
,
.CAHBLTl0II
(
CAHBLTIlll
)
,
.CAHBLTO1II
(
CAHBLTllll
)
,
.CAHBLTI1II
(
CAHBLTO0ll
)
,
.CAHBLTl1II
(
{
CAHBLTIO0OI
,
CAHBLTOllOI
,
CAHBLTl0IOI
,
CAHBLTIOIOI
,
CAHBLTOlOOI
,
CAHBLTl011
,
CAHBLTIO11
,
CAHBLTOl01
,
CAHBLTl0l1
,
CAHBLTIOl1
,
CAHBLTOlI1
,
CAHBLTl0O1
,
CAHBLTIOO1
,
CAHBLTOl10
,
CAHBLTl000
,
CAHBLTIO00
,
CAHBLTOll0
}
)
,
.CAHBLTOOlI
(
{
CAHBLTlO0OI
,
CAHBLTIllOI
,
CAHBLTO1IOI
,
CAHBLTlOIOI
,
CAHBLTIlOOI
,
CAHBLTO111
,
CAHBLTlO11
,
CAHBLTIl01
,
CAHBLTO1l1
,
CAHBLTlOl1
,
CAHBLTIlI1
,
CAHBLTO1O1
,
CAHBLTlOO1
,
CAHBLTIl10
,
CAHBLTO100
,
CAHBLTlO00
,
CAHBLTIll0
}
)
,
.CAHBLTIOlI
(
CAHBLTl0O0
[
15
:
0
]
)
,
.CAHBLTlOlI
(
CAHBLTl00OI
)
,
.CAHBLTOIlI
(
CAHBLTO10OI
)
,
.CAHBLTIIlI
(
CAHBLTlIl0
)
,
.HRDATA_S0
(
CAHBLTllI0I
)
,
.HREADYOUT_S0
(
CAHBLTO100I
)
,
.HRDATA_S1
(
CAHBLTO0I0I
)
,
.HREADYOUT_S1
(
CAHBLTI100I
)
,
.HRDATA_S2
(
CAHBLTI0I0I
)
,
.HREADYOUT_S2
(
CAHBLTl100I
)
,
.HRDATA_S3
(
CAHBLTl0I0I
)
,
.HREADYOUT_S3
(
CAHBLTOO10I
)
,
.HRDATA_S4
(
CAHBLTO1I0I
)
,
.HREADYOUT_S4
(
CAHBLTIO10I
)
,
.HRDATA_S5
(
CAHBLTI1I0I
)
,
.HREADYOUT_S5
(
CAHBLTlO10I
)
,
.HRDATA_S6
(
CAHBLTl1I0I
)
,
.HREADYOUT_S6
(
CAHBLTOI10I
)
,
.HRDATA_S7
(
CAHBLTOOl0I
)
,
.HREADYOUT_S7
(
CAHBLTII10I
)
,
.HRDATA_S8
(
CAHBLTIOl0I
)
,
.HREADYOUT_S8
(
CAHBLTlI10I
)
,
.HRDATA_S9
(
CAHBLTlOl0I
)
,
.HREADYOUT_S9
(
CAHBLTOl10I
)
,
.HRDATA_S10
(
CAHBLTOIl0I
)
,
.HREADYOUT_S10
(
CAHBLTIl10I
)
,
.HRDATA_S11
(
CAHBLTIIl0I
)
,
.HREADYOUT_S11
(
CAHBLTll10I
)
,
.HRDATA_S12
(
CAHBLTlIl0I
)
,
.HREADYOUT_S12
(
CAHBLTO010I
)
,
.HRDATA_S13
(
CAHBLTOll0I
)
,
.HREADYOUT_S13
(
CAHBLTI010I
)
,
.HRDATA_S14
(
CAHBLTIll0I
)
,
.HREADYOUT_S14
(
CAHBLTl010I
)
,
.HRDATA_S15
(
CAHBLTlll0I
)
,
.HREADYOUT_S15
(
CAHBLTO110I
)
,
.HRDATA_SHG
(
CAHBLTO0l0I
)
,
.HREADYOUT_SHG
(
CAHBLTI110I
)
,
.CAHBLTlIlI
(
CAHBLTl110I
)
)
;
CAHBLTO0OI
#
(
.MODE_CFG
(
MODE_CFG
)
,
.CAHBLTI
(
CAHBLTIIl0
)
,
.CAHBLTl
(
CAHBLTI0O0
)
)
CAHBLTIlO0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTII
(
1
'b
0
)
,
.CAHBLTI0OI
(
HADDR_M1
)
,
.CAHBLTl0OI
(
HMASTLOCK_M1
)
,
.CAHBLTO1OI
(
HSIZE_M1
)
,
.CAHBLTI1OI
(
HTRANS_M1
)
,
.CAHBLTl1OI
(
HWRITE_M1
)
,
.CAHBLTOOII
(
HRESP_M1
)
,
.CAHBLTIOII
(
HRDATA_M1
)
,
.CAHBLTlOII
(
CAHBLTlIO0l
)
,
.CAHBLTOIII
(
{
CAHBLTO0O0I
,
CAHBLTl11lI
,
CAHBLTII1lI
,
CAHBLTO00lI
,
CAHBLTl1llI
,
CAHBLTIIllI
,
CAHBLTO0IlI
,
CAHBLTl1OlI
,
CAHBLTIIOlI
,
CAHBLTO01II
,
CAHBLTl10II
,
CAHBLTII0II
,
CAHBLTO0lII
,
CAHBLTl1III
,
CAHBLTIIIII
,
CAHBLTO0OII
,
CAHBLTl11OI
}
)
,
.CAHBLTIIII
(
{
CAHBLTI0O0I
,
CAHBLTOOO0I
,
CAHBLTlI1lI
,
CAHBLTI00lI
,
CAHBLTOO0lI
,
CAHBLTlIllI
,
CAHBLTI0IlI
,
CAHBLTOOIlI
,
CAHBLTlIOlI
,
CAHBLTI01II
,
CAHBLTOO1II
,
CAHBLTlI0II
,
CAHBLTI0lII
,
CAHBLTOOlII
,
CAHBLTlIIII
,
CAHBLTI0OII
,
CAHBLTOOOII
}
)
,
.CAHBLTlIII
(
{
CAHBLTl0O0I
,
CAHBLTIOO0I
,
CAHBLTOl1lI
,
CAHBLTl00lI
,
CAHBLTIO0lI
,
CAHBLTOlllI
,
CAHBLTl0IlI
,
CAHBLTIOIlI
,
CAHBLTOlOlI
,
CAHBLTl01II
,
CAHBLTIO1II
,
CAHBLTOl0II
,
CAHBLTl0lII
,
CAHBLTIOlII
,
CAHBLTOlIII
,
CAHBLTl0OII
,
CAHBLTIOOII
}
)
,
.CAHBLTOlII
(
CAHBLTIII0I
)
,
.CAHBLTIlII
(
CAHBLTlII0I
)
,
.CAHBLTllII
(
CAHBLTOlI0I
)
,
.CAHBLTO0II
(
CAHBLTI0ll
)
,
.CAHBLTI0II
(
CAHBLTO01
)
,
.CAHBLTl0II
(
CAHBLTl0ll
)
,
.CAHBLTO1II
(
CAHBLTO1ll
)
,
.CAHBLTI1II
(
CAHBLTI1ll
)
,
.CAHBLTl1II
(
{
CAHBLTlOO0I
,
CAHBLTIl1lI
,
CAHBLTO10lI
,
CAHBLTlO0lI
,
CAHBLTIlllI
,
CAHBLTO1IlI
,
CAHBLTlOIlI
,
CAHBLTIlOlI
,
CAHBLTO11II
,
CAHBLTlO1II
,
CAHBLTIl0II
,
CAHBLTO1lII
,
CAHBLTlOlII
,
CAHBLTIlIII
,
CAHBLTO1OII
,
CAHBLTlOOII
,
CAHBLTIl1OI
}
)
,
.CAHBLTOOlI
(
{
CAHBLTOIO0I
,
CAHBLTll1lI
,
CAHBLTI10lI
,
CAHBLTOI0lI
,
CAHBLTllllI
,
CAHBLTI1IlI
,
CAHBLTOIIlI
,
CAHBLTllOlI
,
CAHBLTI11II
,
CAHBLTOI1II
,
CAHBLTll0II
,
CAHBLTI1lII
,
CAHBLTOIlII
,
CAHBLTllIII
,
CAHBLTI1OII
,
CAHBLTOIOII
,
CAHBLTll1OI
}
)
,
.CAHBLTIOlI
(
CAHBLTO1O0
[
15
:
0
]
)
,
.CAHBLTlOlI
(
CAHBLTO1O0I
)
,
.CAHBLTOIlI
(
CAHBLTI1O0I
)
,
.CAHBLTIIlI
(
CAHBLTOl1OI
)
,
.HRDATA_S0
(
CAHBLTI0l0I
)
,
.HREADYOUT_S0
(
CAHBLTOOO1I
)
,
.HRDATA_S1
(
CAHBLTl0l0I
)
,
.HREADYOUT_S1
(
CAHBLTIOO1I
)
,
.HRDATA_S2
(
CAHBLTO1l0I
)
,
.HREADYOUT_S2
(
CAHBLTlOO1I
)
,
.HRDATA_S3
(
CAHBLTI1l0I
)
,
.HREADYOUT_S3
(
CAHBLTOIO1I
)
,
.HRDATA_S4
(
CAHBLTl1l0I
)
,
.HREADYOUT_S4
(
CAHBLTIIO1I
)
,
.HRDATA_S5
(
CAHBLTOO00I
)
,
.HREADYOUT_S5
(
CAHBLTlIO1I
)
,
.HRDATA_S6
(
CAHBLTIO00I
)
,
.HREADYOUT_S6
(
CAHBLTOlO1I
)
,
.HRDATA_S7
(
CAHBLTlO00I
)
,
.HREADYOUT_S7
(
CAHBLTIlO1I
)
,
.HRDATA_S8
(
CAHBLTOI00I
)
,
.HREADYOUT_S8
(
CAHBLTllO1I
)
,
.HRDATA_S9
(
CAHBLTII00I
)
,
.HREADYOUT_S9
(
CAHBLTO0O1I
)
,
.HRDATA_S10
(
CAHBLTlI00I
)
,
.HREADYOUT_S10
(
CAHBLTI0O1I
)
,
.HRDATA_S11
(
CAHBLTOl00I
)
,
.HREADYOUT_S11
(
CAHBLTl0O1I
)
,
.HRDATA_S12
(
CAHBLTIl00I
)
,
.HREADYOUT_S12
(
CAHBLTO1O1I
)
,
.HRDATA_S13
(
CAHBLTll00I
)
,
.HREADYOUT_S13
(
CAHBLTI1O1I
)
,
.HRDATA_S14
(
CAHBLTO000I
)
,
.HREADYOUT_S14
(
CAHBLTl1O1I
)
,
.HRDATA_S15
(
CAHBLTI000I
)
,
.HREADYOUT_S15
(
CAHBLTOOI1I
)
,
.HRDATA_SHG
(
CAHBLTl000I
)
,
.HREADYOUT_SHG
(
CAHBLTIOI1I
)
,
.CAHBLTlIlI
(
CAHBLTlOI1I
)
)
;
CAHBLTl0Il
CAHBLTllO0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTOII1I
)
,
.CAHBLTOOII
(
CAHBLTlIl1I
)
,
.CAHBLTI1Il
(
HSEL_S0
)
,
.CAHBLTI0OI
(
HADDR_S0
)
,
.CAHBLTO1OI
(
HSIZE_S0
)
,
.CAHBLTI1OI
(
HTRANS_S0
)
,
.CAHBLTl1OI
(
HWRITE_S0
)
,
.CAHBLTl1Il
(
HWDATA_S0
)
,
.CAHBLTOOll
(
HREADY_S0
)
,
.CAHBLTl0OI
(
HMASTLOCK_S0
)
,
.CAHBLTOl1
(
{
CAHBLTO11OI
,
CAHBLTl0l0
}
)
,
.CAHBLTIOll
(
{
CAHBLTI11OI
,
CAHBLTO1l0
}
)
,
.CAHBLTlOll
(
{
CAHBLTIO1ll
,
CAHBLTI1lll
}
)
,
.CAHBLTOIll
(
{
CAHBLTO01OI
,
CAHBLTlll0
}
)
,
.CAHBLTIIll
(
{
CAHBLTI01OI
,
CAHBLTO0l0
}
)
,
.CAHBLTlIll
(
{
CAHBLTl01OI
,
CAHBLTI0l0
}
)
,
.CAHBLTOlll
(
CAHBLTI1OOl
)
,
.CAHBLTll1
(
CAHBLTI0OIl
)
,
.CAHBLTIlll
(
CAHBLTII0Ol
)
,
.CAHBLTllll
(
CAHBLTIO0Il
)
,
.CAHBLTO0ll
(
CAHBLTIlOll
)
,
.CAHBLTI0ll
(
CAHBLTIOlOl
)
,
.CAHBLTO01
(
CAHBLTI1IIl
)
,
.CAHBLTl0ll
(
CAHBLTIl1Ol
)
,
.CAHBLTO1ll
(
CAHBLTII1Il
)
,
.CAHBLTI1ll
(
CAHBLTI0Ill
)
,
.HWDATA_M0
(
CAHBLTIl01I
)
,
.HWDATA_M1
(
CAHBLTI011I
)
)
;
CAHBLTl0Il
CAHBLTO0O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTIII1I
)
,
.CAHBLTOOII
(
CAHBLTOll1I
)
,
.CAHBLTI1Il
(
HSEL_S1
)
,
.CAHBLTI0OI
(
HADDR_S1
)
,
.CAHBLTO1OI
(
HSIZE_S1
)
,
.CAHBLTI1OI
(
HTRANS_S1
)
,
.CAHBLTl1OI
(
HWRITE_S1
)
,
.CAHBLTl1Il
(
HWDATA_S1
)
,
.CAHBLTOOll
(
HREADY_S1
)
,
.CAHBLTl0OI
(
HMASTLOCK_S1
)
,
.CAHBLTOl1
(
{
CAHBLTIlOII
,
CAHBLTOl00
}
)
,
.CAHBLTIOll
(
{
CAHBLTllOII
,
CAHBLTIl00
}
)
,
.CAHBLTlOll
(
{
CAHBLTlO1ll
,
CAHBLTl1lll
}
)
,
.CAHBLTOIll
(
{
CAHBLTIIOII
,
CAHBLTOI00
}
)
,
.CAHBLTIIll
(
{
CAHBLTlIOII
,
CAHBLTII00
}
)
,
.CAHBLTlIll
(
{
CAHBLTOlOII
,
CAHBLTlI00
}
)
,
.CAHBLTOlll
(
CAHBLTl1OOl
)
,
.CAHBLTll1
(
CAHBLTl0OIl
)
,
.CAHBLTIlll
(
CAHBLTlI0Ol
)
,
.CAHBLTllll
(
CAHBLTlO0Il
)
,
.CAHBLTO0ll
(
CAHBLTllOll
)
,
.CAHBLTI0ll
(
CAHBLTlOlOl
)
,
.CAHBLTO01
(
CAHBLTl1IIl
)
,
.CAHBLTl0ll
(
CAHBLTll1Ol
)
,
.CAHBLTO1ll
(
CAHBLTlI1Il
)
,
.CAHBLTI1ll
(
CAHBLTl0Ill
)
,
.HWDATA_M0
(
CAHBLTll01I
)
,
.HWDATA_M1
(
CAHBLTl011I
)
)
;
CAHBLTl0Il
CAHBLTI0O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTlII1I
)
,
.CAHBLTOOII
(
CAHBLTIll1I
)
,
.CAHBLTI1Il
(
HSEL_S2
)
,
.CAHBLTI0OI
(
HADDR_S2
)
,
.CAHBLTO1OI
(
HSIZE_S2
)
,
.CAHBLTI1OI
(
HTRANS_S2
)
,
.CAHBLTl1OI
(
HWRITE_S2
)
,
.CAHBLTl1Il
(
HWDATA_S2
)
,
.CAHBLTOOll
(
HREADY_S2
)
,
.CAHBLTl0OI
(
HMASTLOCK_S2
)
,
.CAHBLTOl1
(
{
CAHBLTlOIII
,
CAHBLTIO10
}
)
,
.CAHBLTIOll
(
{
CAHBLTOIIII
,
CAHBLTlO10
}
)
,
.CAHBLTlOll
(
{
CAHBLTOI1ll
,
CAHBLTOO0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTl1OII
,
CAHBLTI100
}
)
,
.CAHBLTIIll
(
{
CAHBLTOOIII
,
CAHBLTl100
}
)
,
.CAHBLTlIll
(
{
CAHBLTIOIII
,
CAHBLTOO10
}
)
,
.CAHBLTOlll
(
CAHBLTOOIOl
)
,
.CAHBLTll1
(
CAHBLTO1OIl
)
,
.CAHBLTIlll
(
CAHBLTOl0Ol
)
,
.CAHBLTllll
(
CAHBLTOI0Il
)
,
.CAHBLTO0ll
(
CAHBLTO0Oll
)
,
.CAHBLTI0ll
(
CAHBLTOIlOl
)
,
.CAHBLTO01
(
CAHBLTOOlIl
)
,
.CAHBLTl0ll
(
CAHBLTO01Ol
)
,
.CAHBLTO1ll
(
CAHBLTOl1Il
)
,
.CAHBLTI1ll
(
CAHBLTO1Ill
)
,
.HWDATA_M0
(
CAHBLTO001I
)
,
.HWDATA_M1
(
CAHBLTO111I
)
)
;
CAHBLTl0Il
CAHBLTl0O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTOlI1I
)
,
.CAHBLTOOII
(
CAHBLTlll1I
)
,
.CAHBLTI1Il
(
HSEL_S3
)
,
.CAHBLTI0OI
(
HADDR_S3
)
,
.CAHBLTO1OI
(
HSIZE_S3
)
,
.CAHBLTI1OI
(
HTRANS_S3
)
,
.CAHBLTl1OI
(
HWRITE_S3
)
,
.CAHBLTl1Il
(
HWDATA_S3
)
,
.CAHBLTOOll
(
HREADY_S3
)
,
.CAHBLTl0OI
(
HMASTLOCK_S3
)
,
.CAHBLTOl1
(
{
CAHBLTO1III
,
CAHBLTl010
}
)
,
.CAHBLTIOll
(
{
CAHBLTI1III
,
CAHBLTO110
}
)
,
.CAHBLTlOll
(
{
CAHBLTII1ll
,
CAHBLTIO0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTO0III
,
CAHBLTll10
}
)
,
.CAHBLTIIll
(
{
CAHBLTI0III
,
CAHBLTO010
}
)
,
.CAHBLTlIll
(
{
CAHBLTl0III
,
CAHBLTI010
}
)
,
.CAHBLTOlll
(
CAHBLTIOIOl
)
,
.CAHBLTll1
(
CAHBLTI1OIl
)
,
.CAHBLTIlll
(
CAHBLTIl0Ol
)
,
.CAHBLTllll
(
CAHBLTII0Il
)
,
.CAHBLTO0ll
(
CAHBLTI0Oll
)
,
.CAHBLTI0ll
(
CAHBLTIIlOl
)
,
.CAHBLTO01
(
CAHBLTIOlIl
)
,
.CAHBLTl0ll
(
CAHBLTI01Ol
)
,
.CAHBLTO1ll
(
CAHBLTIl1Il
)
,
.CAHBLTI1ll
(
CAHBLTI1Ill
)
,
.HWDATA_M0
(
CAHBLTI001I
)
,
.HWDATA_M1
(
CAHBLTI111I
)
)
;
CAHBLTl0Il
CAHBLTO1O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTIlI1I
)
,
.CAHBLTOOII
(
CAHBLTO0l1I
)
,
.CAHBLTI1Il
(
HSEL_S4
)
,
.CAHBLTI0OI
(
HADDR_S4
)
,
.CAHBLTO1OI
(
HSIZE_S4
)
,
.CAHBLTI1OI
(
HTRANS_S4
)
,
.CAHBLTl1OI
(
HWRITE_S4
)
,
.CAHBLTl1Il
(
HWDATA_S4
)
,
.CAHBLTOOll
(
HREADY_S4
)
,
.CAHBLTl0OI
(
HMASTLOCK_S4
)
,
.CAHBLTOl1
(
{
CAHBLTIllII
,
CAHBLTOlO1
}
)
,
.CAHBLTIOll
(
{
CAHBLTlllII
,
CAHBLTIlO1
}
)
,
.CAHBLTlOll
(
{
CAHBLTlI1ll
,
CAHBLTlO0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTIIlII
,
CAHBLTOIO1
}
)
,
.CAHBLTIIll
(
{
CAHBLTlIlII
,
CAHBLTIIO1
}
)
,
.CAHBLTlIll
(
{
CAHBLTOllII
,
CAHBLTlIO1
}
)
,
.CAHBLTOlll
(
CAHBLTlOIOl
)
,
.CAHBLTll1
(
CAHBLTl1OIl
)
,
.CAHBLTIlll
(
CAHBLTll0Ol
)
,
.CAHBLTllll
(
CAHBLTlI0Il
)
,
.CAHBLTO0ll
(
CAHBLTl0Oll
)
,
.CAHBLTI0ll
(
CAHBLTlIlOl
)
,
.CAHBLTO01
(
CAHBLTlOlIl
)
,
.CAHBLTl0ll
(
CAHBLTl01Ol
)
,
.CAHBLTO1ll
(
CAHBLTll1Il
)
,
.CAHBLTI1ll
(
CAHBLTl1Ill
)
,
.HWDATA_M0
(
CAHBLTl001I
)
,
.HWDATA_M1
(
CAHBLTl111I
)
)
;
CAHBLTl0Il
CAHBLTI1O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTllI1I
)
,
.CAHBLTOOII
(
CAHBLTI0l1I
)
,
.CAHBLTI1Il
(
HSEL_S5
)
,
.CAHBLTI0OI
(
HADDR_S5
)
,
.CAHBLTO1OI
(
HSIZE_S5
)
,
.CAHBLTI1OI
(
HTRANS_S5
)
,
.CAHBLTl1OI
(
HWRITE_S5
)
,
.CAHBLTl1Il
(
HWDATA_S5
)
,
.CAHBLTOOll
(
HREADY_S5
)
,
.CAHBLTl0OI
(
HMASTLOCK_S5
)
,
.CAHBLTOl1
(
{
CAHBLTlO0II
,
CAHBLTIOI1
}
)
,
.CAHBLTIOll
(
{
CAHBLTOI0II
,
CAHBLTlOI1
}
)
,
.CAHBLTlOll
(
{
CAHBLTOl1ll
,
CAHBLTOI0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTl1lII
,
CAHBLTI1O1
}
)
,
.CAHBLTIIll
(
{
CAHBLTOO0II
,
CAHBLTl1O1
}
)
,
.CAHBLTlIll
(
{
CAHBLTIO0II
,
CAHBLTOOI1
}
)
,
.CAHBLTOlll
(
CAHBLTOIIOl
)
,
.CAHBLTll1
(
CAHBLTOOIIl
)
,
.CAHBLTIlll
(
CAHBLTO00Ol
)
,
.CAHBLTllll
(
CAHBLTOl0Il
)
,
.CAHBLTO0ll
(
CAHBLTO1Oll
)
,
.CAHBLTI0ll
(
CAHBLTOllOl
)
,
.CAHBLTO01
(
CAHBLTOIlIl
)
,
.CAHBLTl0ll
(
CAHBLTO11Ol
)
,
.CAHBLTO1ll
(
CAHBLTO01Il
)
,
.CAHBLTI1ll
(
CAHBLTOOlll
)
,
.HWDATA_M0
(
CAHBLTO101I
)
,
.HWDATA_M1
(
CAHBLTOOOOl
)
)
;
CAHBLTl0Il
CAHBLTl1O0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTO0I1I
)
,
.CAHBLTOOII
(
CAHBLTl0l1I
)
,
.CAHBLTI1Il
(
HSEL_S6
)
,
.CAHBLTI0OI
(
HADDR_S6
)
,
.CAHBLTO1OI
(
HSIZE_S6
)
,
.CAHBLTI1OI
(
HTRANS_S6
)
,
.CAHBLTl1OI
(
HWRITE_S6
)
,
.CAHBLTl1Il
(
HWDATA_S6
)
,
.CAHBLTOOll
(
HREADY_S6
)
,
.CAHBLTl0OI
(
HMASTLOCK_S6
)
,
.CAHBLTOl1
(
{
CAHBLTO10II
,
CAHBLTl0I1
}
)
,
.CAHBLTIOll
(
{
CAHBLTI10II
,
CAHBLTO1I1
}
)
,
.CAHBLTlOll
(
{
CAHBLTIl1ll
,
CAHBLTII0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTO00II
,
CAHBLTllI1
}
)
,
.CAHBLTIIll
(
{
CAHBLTI00II
,
CAHBLTO0I1
}
)
,
.CAHBLTlIll
(
{
CAHBLTl00II
,
CAHBLTI0I1
}
)
,
.CAHBLTOlll
(
CAHBLTIIIOl
)
,
.CAHBLTll1
(
CAHBLTIOIIl
)
,
.CAHBLTIlll
(
CAHBLTI00Ol
)
,
.CAHBLTllll
(
CAHBLTIl0Il
)
,
.CAHBLTO0ll
(
CAHBLTI1Oll
)
,
.CAHBLTI0ll
(
CAHBLTIllOl
)
,
.CAHBLTO01
(
CAHBLTIIlIl
)
,
.CAHBLTl0ll
(
CAHBLTI11Ol
)
,
.CAHBLTO1ll
(
CAHBLTI01Il
)
,
.CAHBLTI1ll
(
CAHBLTIOlll
)
,
.HWDATA_M0
(
CAHBLTI101I
)
,
.HWDATA_M1
(
CAHBLTIOOOl
)
)
;
CAHBLTl0Il
CAHBLTOOI0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTI0I1I
)
,
.CAHBLTOOII
(
CAHBLTO1l1I
)
,
.CAHBLTI1Il
(
HSEL_S7
)
,
.CAHBLTI0OI
(
HADDR_S7
)
,
.CAHBLTO1OI
(
HSIZE_S7
)
,
.CAHBLTI1OI
(
HTRANS_S7
)
,
.CAHBLTl1OI
(
HWRITE_S7
)
,
.CAHBLTl1Il
(
HWDATA_S7
)
,
.CAHBLTOOll
(
HREADY_S7
)
,
.CAHBLTl0OI
(
HMASTLOCK_S7
)
,
.CAHBLTOl1
(
{
CAHBLTIl1II
,
CAHBLTOll1
}
)
,
.CAHBLTIOll
(
{
CAHBLTll1II
,
CAHBLTIll1
}
)
,
.CAHBLTlOll
(
{
CAHBLTll1ll
,
CAHBLTlI0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTII1II
,
CAHBLTOIl1
}
)
,
.CAHBLTIIll
(
{
CAHBLTlI1II
,
CAHBLTIIl1
}
)
,
.CAHBLTlIll
(
{
CAHBLTOl1II
,
CAHBLTlIl1
}
)
,
.CAHBLTOlll
(
CAHBLTlIIOl
)
,
.CAHBLTll1
(
CAHBLTlOIIl
)
,
.CAHBLTIlll
(
CAHBLTl00Ol
)
,
.CAHBLTllll
(
CAHBLTll0Il
)
,
.CAHBLTO0ll
(
CAHBLTl1Oll
)
,
.CAHBLTI0ll
(
CAHBLTlllOl
)
,
.CAHBLTO01
(
CAHBLTlIlIl
)
,
.CAHBLTl0ll
(
CAHBLTl11Ol
)
,
.CAHBLTO1ll
(
CAHBLTl01Il
)
,
.CAHBLTI1ll
(
CAHBLTlOlll
)
,
.HWDATA_M0
(
CAHBLTl101I
)
,
.HWDATA_M1
(
CAHBLTlOOOl
)
)
;
CAHBLTl0Il
CAHBLTIOI0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTl0I1I
)
,
.CAHBLTOOII
(
CAHBLTI1l1I
)
,
.CAHBLTI1Il
(
HSEL_S8
)
,
.CAHBLTI0OI
(
HADDR_S8
)
,
.CAHBLTO1OI
(
HSIZE_S8
)
,
.CAHBLTI1OI
(
HTRANS_S8
)
,
.CAHBLTl1OI
(
HWRITE_S8
)
,
.CAHBLTl1Il
(
HWDATA_S8
)
,
.CAHBLTOOll
(
HREADY_S8
)
,
.CAHBLTl0OI
(
HMASTLOCK_S8
)
,
.CAHBLTOl1
(
{
CAHBLTlOOlI
,
CAHBLTIO01
}
)
,
.CAHBLTIOll
(
{
CAHBLTOIOlI
,
CAHBLTlO01
}
)
,
.CAHBLTlOll
(
{
CAHBLTO01ll
,
CAHBLTOl0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTl11II
,
CAHBLTI1l1
}
)
,
.CAHBLTIIll
(
{
CAHBLTOOOlI
,
CAHBLTl1l1
}
)
,
.CAHBLTlIll
(
{
CAHBLTIOOlI
,
CAHBLTOO01
}
)
,
.CAHBLTOlll
(
CAHBLTOlIOl
)
,
.CAHBLTll1
(
CAHBLTOIIIl
)
,
.CAHBLTIlll
(
CAHBLTO10Ol
)
,
.CAHBLTllll
(
CAHBLTO00Il
)
,
.CAHBLTO0ll
(
CAHBLTOOIll
)
,
.CAHBLTI0ll
(
CAHBLTO0lOl
)
,
.CAHBLTO01
(
CAHBLTOllIl
)
,
.CAHBLTl0ll
(
CAHBLTOOOIl
)
,
.CAHBLTO1ll
(
CAHBLTO11Il
)
,
.CAHBLTI1ll
(
CAHBLTOIlll
)
,
.HWDATA_M0
(
CAHBLTOO11I
)
,
.HWDATA_M1
(
CAHBLTOIOOl
)
)
;
CAHBLTl0Il
CAHBLTlOI0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTO1I1I
)
,
.CAHBLTOOII
(
CAHBLTl1l1I
)
,
.CAHBLTI1Il
(
HSEL_S9
)
,
.CAHBLTI0OI
(
HADDR_S9
)
,
.CAHBLTO1OI
(
HSIZE_S9
)
,
.CAHBLTI1OI
(
HTRANS_S9
)
,
.CAHBLTl1OI
(
HWRITE_S9
)
,
.CAHBLTl1Il
(
HWDATA_S9
)
,
.CAHBLTOOll
(
HREADY_S9
)
,
.CAHBLTl0OI
(
HMASTLOCK_S9
)
,
.CAHBLTOl1
(
{
CAHBLTO1OlI
,
CAHBLTl001
}
)
,
.CAHBLTIOll
(
{
CAHBLTI1OlI
,
CAHBLTO101
}
)
,
.CAHBLTlOll
(
{
CAHBLTI01ll
,
CAHBLTIl0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTO0OlI
,
CAHBLTll01
}
)
,
.CAHBLTIIll
(
{
CAHBLTI0OlI
,
CAHBLTO001
}
)
,
.CAHBLTlIll
(
{
CAHBLTl0OlI
,
CAHBLTI001
}
)
,
.CAHBLTOlll
(
CAHBLTIlIOl
)
,
.CAHBLTll1
(
CAHBLTIIIIl
)
,
.CAHBLTIlll
(
CAHBLTI10Ol
)
,
.CAHBLTllll
(
CAHBLTI00Il
)
,
.CAHBLTO0ll
(
CAHBLTIOIll
)
,
.CAHBLTI0ll
(
CAHBLTI0lOl
)
,
.CAHBLTO01
(
CAHBLTIllIl
)
,
.CAHBLTl0ll
(
CAHBLTIOOIl
)
,
.CAHBLTO1ll
(
CAHBLTI11Il
)
,
.CAHBLTI1ll
(
CAHBLTIIlll
)
,
.HWDATA_M0
(
CAHBLTIO11I
)
,
.HWDATA_M1
(
CAHBLTIIOOl
)
)
;
CAHBLTl0Il
CAHBLTOII0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTI1I1I
)
,
.CAHBLTOOII
(
CAHBLTOO01I
)
,
.CAHBLTI1Il
(
HSEL_S10
)
,
.CAHBLTI0OI
(
HADDR_S10
)
,
.CAHBLTO1OI
(
HSIZE_S10
)
,
.CAHBLTI1OI
(
HTRANS_S10
)
,
.CAHBLTl1OI
(
HWRITE_S10
)
,
.CAHBLTl1Il
(
HWDATA_S10
)
,
.CAHBLTOOll
(
HREADY_S10
)
,
.CAHBLTl0OI
(
HMASTLOCK_S10
)
,
.CAHBLTOl1
(
{
CAHBLTIlIlI
,
CAHBLTOl11
}
)
,
.CAHBLTIOll
(
{
CAHBLTllIlI
,
CAHBLTIl11
}
)
,
.CAHBLTlOll
(
{
CAHBLTl01ll
,
CAHBLTll0ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTIIIlI
,
CAHBLTOI11
}
)
,
.CAHBLTIIll
(
{
CAHBLTlIIlI
,
CAHBLTII11
}
)
,
.CAHBLTlIll
(
{
CAHBLTOlIlI
,
CAHBLTlI11
}
)
,
.CAHBLTOlll
(
CAHBLTllIOl
)
,
.CAHBLTll1
(
CAHBLTlIIIl
)
,
.CAHBLTIlll
(
CAHBLTl10Ol
)
,
.CAHBLTllll
(
CAHBLTl00Il
)
,
.CAHBLTO0ll
(
CAHBLTlOIll
)
,
.CAHBLTI0ll
(
CAHBLTl0lOl
)
,
.CAHBLTO01
(
CAHBLTlllIl
)
,
.CAHBLTl0ll
(
CAHBLTlOOIl
)
,
.CAHBLTO1ll
(
CAHBLTl11Il
)
,
.CAHBLTI1ll
(
CAHBLTlIlll
)
,
.HWDATA_M0
(
CAHBLTlO11I
)
,
.HWDATA_M1
(
CAHBLTlIOOl
)
)
;
CAHBLTl0Il
CAHBLTIII0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTl1I1I
)
,
.CAHBLTOOII
(
CAHBLTIO01I
)
,
.CAHBLTI1Il
(
HSEL_S11
)
,
.CAHBLTI0OI
(
HADDR_S11
)
,
.CAHBLTO1OI
(
HSIZE_S11
)
,
.CAHBLTI1OI
(
HTRANS_S11
)
,
.CAHBLTl1OI
(
HWRITE_S11
)
,
.CAHBLTl1Il
(
HWDATA_S11
)
,
.CAHBLTOOll
(
HREADY_S11
)
,
.CAHBLTl0OI
(
HMASTLOCK_S11
)
,
.CAHBLTOl1
(
{
CAHBLTlOllI
,
CAHBLTIOOOI
}
)
,
.CAHBLTIOll
(
{
CAHBLTOIllI
,
CAHBLTlOOOI
}
)
,
.CAHBLTlOll
(
{
CAHBLTO11ll
,
CAHBLTO00ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTl1IlI
,
CAHBLTI111
}
)
,
.CAHBLTIIll
(
{
CAHBLTOOllI
,
CAHBLTl111
}
)
,
.CAHBLTlIll
(
{
CAHBLTIOllI
,
CAHBLTOOOOI
}
)
,
.CAHBLTOlll
(
CAHBLTO0IOl
)
,
.CAHBLTll1
(
CAHBLTOlIIl
)
,
.CAHBLTIlll
(
CAHBLTOO1Ol
)
,
.CAHBLTllll
(
CAHBLTO10Il
)
,
.CAHBLTO0ll
(
CAHBLTOIIll
)
,
.CAHBLTI0ll
(
CAHBLTO1lOl
)
,
.CAHBLTO01
(
CAHBLTO0lIl
)
,
.CAHBLTl0ll
(
CAHBLTOIOIl
)
,
.CAHBLTO1ll
(
CAHBLTOOOll
)
,
.CAHBLTI1ll
(
CAHBLTOllll
)
,
.HWDATA_M0
(
CAHBLTOI11I
)
,
.HWDATA_M1
(
CAHBLTOlOOl
)
)
;
CAHBLTl0Il
CAHBLTlII0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTOOl1I
)
,
.CAHBLTOOII
(
CAHBLTlO01I
)
,
.CAHBLTI1Il
(
HSEL_S12
)
,
.CAHBLTI0OI
(
HADDR_S12
)
,
.CAHBLTO1OI
(
HSIZE_S12
)
,
.CAHBLTI1OI
(
HTRANS_S12
)
,
.CAHBLTl1OI
(
HWRITE_S12
)
,
.CAHBLTl1Il
(
HWDATA_S12
)
,
.CAHBLTOOll
(
HREADY_S12
)
,
.CAHBLTl0OI
(
HMASTLOCK_S12
)
,
.CAHBLTOl1
(
{
CAHBLTO1llI
,
CAHBLTl0OOI
}
)
,
.CAHBLTIOll
(
{
CAHBLTI1llI
,
CAHBLTO1OOI
}
)
,
.CAHBLTlOll
(
{
CAHBLTI11ll
,
CAHBLTI00ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTO0llI
,
CAHBLTllOOI
}
)
,
.CAHBLTIIll
(
{
CAHBLTI0llI
,
CAHBLTO0OOI
}
)
,
.CAHBLTlIll
(
{
CAHBLTl0llI
,
CAHBLTI0OOI
}
)
,
.CAHBLTOlll
(
CAHBLTI0IOl
)
,
.CAHBLTll1
(
CAHBLTIlIIl
)
,
.CAHBLTIlll
(
CAHBLTIO1Ol
)
,
.CAHBLTllll
(
CAHBLTI10Il
)
,
.CAHBLTO0ll
(
CAHBLTIIIll
)
,
.CAHBLTI0ll
(
CAHBLTI1lOl
)
,
.CAHBLTO01
(
CAHBLTI0lIl
)
,
.CAHBLTl0ll
(
CAHBLTIIOIl
)
,
.CAHBLTO1ll
(
CAHBLTIOOll
)
,
.CAHBLTI1ll
(
CAHBLTIllll
)
,
.HWDATA_M0
(
CAHBLTII11I
)
,
.HWDATA_M1
(
CAHBLTIlOOl
)
)
;
CAHBLTl0Il
CAHBLTOlI0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTIOl1I
)
,
.CAHBLTOOII
(
CAHBLTOI01I
)
,
.CAHBLTI1Il
(
HSEL_S13
)
,
.CAHBLTI0OI
(
HADDR_S13
)
,
.CAHBLTO1OI
(
HSIZE_S13
)
,
.CAHBLTI1OI
(
HTRANS_S13
)
,
.CAHBLTl1OI
(
HWRITE_S13
)
,
.CAHBLTl1Il
(
HWDATA_S13
)
,
.CAHBLTOOll
(
HREADY_S13
)
,
.CAHBLTl0OI
(
HMASTLOCK_S13
)
,
.CAHBLTOl1
(
{
CAHBLTIl0lI
,
CAHBLTOlIOI
}
)
,
.CAHBLTIOll
(
{
CAHBLTll0lI
,
CAHBLTIlIOI
}
)
,
.CAHBLTlOll
(
{
CAHBLTl11ll
,
CAHBLTl00ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTII0lI
,
CAHBLTOIIOI
}
)
,
.CAHBLTIIll
(
{
CAHBLTlI0lI
,
CAHBLTIIIOI
}
)
,
.CAHBLTlIll
(
{
CAHBLTOl0lI
,
CAHBLTlIIOI
}
)
,
.CAHBLTOlll
(
CAHBLTl0IOl
)
,
.CAHBLTll1
(
CAHBLTllIIl
)
,
.CAHBLTIlll
(
CAHBLTlO1Ol
)
,
.CAHBLTllll
(
CAHBLTl10Il
)
,
.CAHBLTO0ll
(
CAHBLTlIIll
)
,
.CAHBLTI0ll
(
CAHBLTl1lOl
)
,
.CAHBLTO01
(
CAHBLTl0lIl
)
,
.CAHBLTl0ll
(
CAHBLTlIOIl
)
,
.CAHBLTO1ll
(
CAHBLTlOOll
)
,
.CAHBLTI1ll
(
CAHBLTlllll
)
,
.HWDATA_M0
(
CAHBLTlI11I
)
,
.HWDATA_M1
(
CAHBLTllOOl
)
)
;
CAHBLTl0Il
CAHBLTIlI0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTlOl1I
)
,
.CAHBLTOOII
(
CAHBLTII01I
)
,
.CAHBLTI1Il
(
HSEL_S14
)
,
.CAHBLTI0OI
(
HADDR_S14
)
,
.CAHBLTO1OI
(
HSIZE_S14
)
,
.CAHBLTI1OI
(
HTRANS_S14
)
,
.CAHBLTl1OI
(
HWRITE_S14
)
,
.CAHBLTl1Il
(
HWDATA_S14
)
,
.CAHBLTOOll
(
HREADY_S14
)
,
.CAHBLTl0OI
(
HMASTLOCK_S14
)
,
.CAHBLTOl1
(
{
CAHBLTlO1lI
,
CAHBLTIOlOI
}
)
,
.CAHBLTIOll
(
{
CAHBLTOI1lI
,
CAHBLTlOlOI
}
)
,
.CAHBLTlOll
(
{
CAHBLTOOO0l
,
CAHBLTO10ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTl10lI
,
CAHBLTI1IOI
}
)
,
.CAHBLTIIll
(
{
CAHBLTOO1lI
,
CAHBLTl1IOI
}
)
,
.CAHBLTlIll
(
{
CAHBLTIO1lI
,
CAHBLTOOlOI
}
)
,
.CAHBLTOlll
(
CAHBLTO1IOl
)
,
.CAHBLTll1
(
CAHBLTO0IIl
)
,
.CAHBLTIlll
(
CAHBLTOI1Ol
)
,
.CAHBLTllll
(
CAHBLTOO1Il
)
,
.CAHBLTO0ll
(
CAHBLTOlIll
)
,
.CAHBLTI0ll
(
CAHBLTOO0Ol
)
,
.CAHBLTO01
(
CAHBLTO1lIl
)
,
.CAHBLTl0ll
(
CAHBLTOlOIl
)
,
.CAHBLTO1ll
(
CAHBLTOIOll
)
,
.CAHBLTI1ll
(
CAHBLTO0lll
)
,
.HWDATA_M0
(
CAHBLTOl11I
)
,
.HWDATA_M1
(
CAHBLTO0OOl
)
)
;
CAHBLTl0Il
CAHBLTllI0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTOIl1I
)
,
.CAHBLTOOII
(
CAHBLTlI01I
)
,
.CAHBLTI1Il
(
HSEL_S15
)
,
.CAHBLTI0OI
(
HADDR_S15
)
,
.CAHBLTO1OI
(
HSIZE_S15
)
,
.CAHBLTI1OI
(
HTRANS_S15
)
,
.CAHBLTl1OI
(
HWRITE_S15
)
,
.CAHBLTl1Il
(
HWDATA_S15
)
,
.CAHBLTOOll
(
HREADY_S15
)
,
.CAHBLTl0OI
(
HMASTLOCK_S15
)
,
.CAHBLTOl1
(
{
CAHBLTO11lI
,
CAHBLTl0lOI
}
)
,
.CAHBLTIOll
(
{
CAHBLTI11lI
,
CAHBLTO1lOI
}
)
,
.CAHBLTlOll
(
{
CAHBLTIOO0l
,
CAHBLTI10ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTO01lI
,
CAHBLTlllOI
}
)
,
.CAHBLTIIll
(
{
CAHBLTI01lI
,
CAHBLTO0lOI
}
)
,
.CAHBLTlIll
(
{
CAHBLTl01lI
,
CAHBLTI0lOI
}
)
,
.CAHBLTOlll
(
CAHBLTI1IOl
)
,
.CAHBLTll1
(
CAHBLTI0IIl
)
,
.CAHBLTIlll
(
CAHBLTII1Ol
)
,
.CAHBLTllll
(
CAHBLTIO1Il
)
,
.CAHBLTO0ll
(
CAHBLTIlIll
)
,
.CAHBLTI0ll
(
CAHBLTIO0Ol
)
,
.CAHBLTO01
(
CAHBLTI1lIl
)
,
.CAHBLTl0ll
(
CAHBLTIlOIl
)
,
.CAHBLTO1ll
(
CAHBLTIIOll
)
,
.CAHBLTI1ll
(
CAHBLTI0lll
)
,
.HWDATA_M0
(
CAHBLTIl11I
)
,
.HWDATA_M1
(
CAHBLTI0OOl
)
)
;
CAHBLTl0Il
CAHBLTO0I0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTIIl1I
)
,
.CAHBLTOOII
(
CAHBLTOl01I
)
,
.CAHBLTI1Il
(
HSEL_SHG
)
,
.CAHBLTI0OI
(
HADDR_SHG
)
,
.CAHBLTO1OI
(
HSIZE_SHG
)
,
.CAHBLTI1OI
(
HTRANS_SHG
)
,
.CAHBLTl1OI
(
HWRITE_SHG
)
,
.CAHBLTl1Il
(
HWDATA_SHG
)
,
.CAHBLTOOll
(
HREADY_SHG
)
,
.CAHBLTl0OI
(
HMASTLOCK_SHG
)
,
.CAHBLTOl1
(
{
CAHBLTIlO0I
,
CAHBLTOl0OI
}
)
,
.CAHBLTIOll
(
{
CAHBLTllO0I
,
CAHBLTIl0OI
}
)
,
.CAHBLTlOll
(
{
CAHBLTlOO0l
,
CAHBLTl10ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTIIO0I
,
CAHBLTOI0OI
}
)
,
.CAHBLTIIll
(
{
CAHBLTlIO0I
,
CAHBLTII0OI
}
)
,
.CAHBLTlIll
(
{
CAHBLTOlO0I
,
CAHBLTlI0OI
}
)
,
.CAHBLTOlll
(
CAHBLTl1IOl
)
,
.CAHBLTll1
(
CAHBLTl0IIl
)
,
.CAHBLTIlll
(
CAHBLTlI1Ol
)
,
.CAHBLTllll
(
CAHBLTlO1Il
)
,
.CAHBLTO0ll
(
CAHBLTllIll
)
,
.CAHBLTI0ll
(
CAHBLTlO0Ol
)
,
.CAHBLTO01
(
CAHBLTl1lIl
)
,
.CAHBLTl0ll
(
CAHBLTllOIl
)
,
.CAHBLTO1ll
(
CAHBLTlIOll
)
,
.CAHBLTI1ll
(
CAHBLTl0lll
)
,
.HWDATA_M0
(
CAHBLTll11I
)
,
.HWDATA_M1
(
CAHBLTl0OOl
)
)
;
CAHBLTllO0
#
(
.MODE_CFG
(
MODE_CFG
)
,
.CAHBLTO0O0
(
CAHBLTO0O0
)
,
.CAHBLTI0O0
(
CAHBLTI0O0
)
)
CAHBLTI0I0l
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTO1Il
(
CAHBLTIlI0I
)
,
.CAHBLTl0O0
(
CAHBLTl0O0
)
,
.CAHBLTO1O0
(
CAHBLTO1O0
)
,
.CAHBLTOl1
(
{
CAHBLTlOI0I
,
CAHBLTIO1OI
}
)
,
.CAHBLTIOll
(
{
CAHBLTOII0I
,
CAHBLTlO1OI
}
)
,
.CAHBLTlOll
(
{
CAHBLTOIO0l
,
CAHBLTOO1ll
}
)
,
.CAHBLTOIll
(
{
CAHBLTl1O0I
,
CAHBLTI10OI
}
)
,
.CAHBLTIIll
(
{
CAHBLTOOI0I
,
CAHBLTl10OI
}
)
,
.CAHBLTlIll
(
{
CAHBLTIOI0I
,
CAHBLTOO1OI
}
)
,
.CAHBLTOlll
(
CAHBLTOOlOl
)
,
.CAHBLTll1
(
CAHBLTO1IIl
)
,
.CAHBLTIlll
(
CAHBLTOl1Ol
)
,
.CAHBLTllll
(
CAHBLTOI1Il
)
,
.CAHBLTO0ll
(
CAHBLTO0Ill
)
,
.CAHBLTI0ll
(
CAHBLTOI0Ol
)
,
.CAHBLTO01
(
CAHBLTOO0Il
)
,
.CAHBLTl0ll
(
CAHBLTO0OIl
)
,
.CAHBLTO1ll
(
CAHBLTOlOll
)
,
.CAHBLTI1ll
(
CAHBLTO1lll
)
,
.HWDATA_M0
(
CAHBLTO011I
)
,
.HWDATA_M1
(
CAHBLTO1OOl
)
,
.CAHBLTll0l
(
CAHBLTll0l
)
,
.CAHBLTO00l
(
CAHBLTO00l
)
,
.CAHBLTI00l
(
CAHBLTI00l
)
,
.CAHBLTl00l
(
CAHBLTl00l
)
)
;
assign
HREADY_M0
=
CAHBLTIIO0l
;
assign
HREADY_M1
=
CAHBLTlIO0l
;
endmodule
