// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 10Feb10		Production Release Version 3.1
// SVN Revision Information:
// SVN $Revision: 11955 $
// SVN $Date: 2010-01-30 15:35:13 -0800 (Sat, 30 Jan 2010) $
`timescale 1ns/1ps
module
CAHBLTlI1
(
input
HCLK,
input
HRESETN,
input
[
1
:
0
]
CAHBLTOl1,
input
CAHBLTIl1,
input
CAHBLTll1,
input
CAHBLTO01,
output
reg
[
1
:
0
]
CAHBLTI01
)
;
localparam
CAHBLTl01
=
3
'b
000
;
localparam
CAHBLTO11
=
3
'b
001
;
localparam
CAHBLTI11
=
3
'b
010
;
localparam
CAHBLTl11
=
3
'b
011
;
localparam
CAHBLTOOOI
=
3
'b
100
;
localparam
CAHBLTIOOI
=
3
'b
101
;
localparam
CAHBLTlOOI
=
3
'b
110
;
localparam
CAHBLTOIOI
=
3
'b
111
;
localparam
CAHBLTIIOI
=
2
'b
01
;
localparam
CAHBLTlIOI
=
2
'b
10
;
localparam
CAHBLTOlOI
=
2
'b
00
;
reg
[
2
:
0
]
CAHBLTIlOI
;
reg
[
2
:
0
]
CAHBLTllOI
;
always
@(*)
begin
CAHBLTI01
=
CAHBLTOlOI
;
case
(
CAHBLTllOI
)
CAHBLTl01
:
begin
if
(
CAHBLTOl1
[
0
]
)
begin
if
(
CAHBLTll1
)
CAHBLTIlOI
=
CAHBLTOOOI
;
else
begin
CAHBLTI01
=
CAHBLTIIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTl11
;
else
CAHBLTIlOI
=
CAHBLTO11
;
end
end
else
if
(
CAHBLTOl1
[
1
]
)
begin
if
(
CAHBLTO01
)
CAHBLTIlOI
=
CAHBLTIOOI
;
else
begin
CAHBLTI01
=
CAHBLTlIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTl01
;
else
CAHBLTIlOI
=
CAHBLTI11
;
end
end
else
CAHBLTIlOI
=
CAHBLTl01
;
end
CAHBLTl11
:
begin
if
(
CAHBLTOl1
[
1
]
)
begin
if
(
CAHBLTO01
)
CAHBLTIlOI
=
CAHBLTIOOI
;
else
begin
CAHBLTI01
=
CAHBLTlIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTl01
;
else
CAHBLTIlOI
=
CAHBLTI11
;
end
end
else
if
(
CAHBLTOl1
[
0
]
)
begin
if
(
CAHBLTll1
)
CAHBLTIlOI
=
CAHBLTOOOI
;
else
begin
CAHBLTI01
=
CAHBLTIIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTl11
;
else
CAHBLTIlOI
=
CAHBLTO11
;
end
end
else
CAHBLTIlOI
=
CAHBLTl11
;
end
CAHBLTO11
:
begin
CAHBLTI01
=
CAHBLTIIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTl11
;
else
CAHBLTIlOI
=
CAHBLTO11
;
end
CAHBLTI11
:
begin
CAHBLTI01
=
CAHBLTlIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTl01
;
else
CAHBLTIlOI
=
CAHBLTI11
;
end
CAHBLTOOOI
:
begin
if
(
CAHBLTll1
)
if
(
CAHBLTOl1
[
0
]
)
begin
CAHBLTI01
=
CAHBLTIIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTOOOI
;
else
CAHBLTIlOI
=
CAHBLTlOOI
;
end
else
CAHBLTIlOI
=
CAHBLTOOOI
;
else
CAHBLTIlOI
=
CAHBLTl11
;
end
CAHBLTlOOI
:
begin
CAHBLTI01
=
CAHBLTIIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTOOOI
;
else
CAHBLTIlOI
=
CAHBLTlOOI
;
end
CAHBLTIOOI
:
begin
if
(
CAHBLTO01
)
if
(
CAHBLTOl1
[
1
]
)
begin
CAHBLTI01
=
CAHBLTlIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTIOOI
;
else
CAHBLTIlOI
=
CAHBLTOIOI
;
end
else
CAHBLTIlOI
=
CAHBLTIOOI
;
else
CAHBLTIlOI
=
CAHBLTl01
;
end
CAHBLTOIOI
:
begin
CAHBLTI01
=
CAHBLTlIOI
;
if
(
CAHBLTIl1
)
CAHBLTIlOI
=
CAHBLTIOOI
;
else
CAHBLTIlOI
=
CAHBLTOIOI
;
end
default
:
CAHBLTIlOI
=
CAHBLTl01
;
endcase
end
always
@
(
posedge
HCLK
or
negedge
HRESETN
)
begin
if
(
!
HRESETN
)
CAHBLTllOI
<=
CAHBLTl01
;
else
CAHBLTllOI
<=
CAHBLTIlOI
;
end
endmodule
