// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 10Feb10		Production Release Version 3.1
// SVN Revision Information:
// SVN $Revision: 11955 $
// SVN $Date: 2010-01-30 15:35:13 -0800 (Sat, 30 Jan 2010) $
`timescale 1ns/1ps
module
CAHBLTO
#
(
parameter
[
0
:
0
]
MODE_CFG
=
0
,
parameter
[
16
:
0
]
CAHBLTI
=
(
2
**
17
)
-
1
,
parameter
[
15
:
0
]
CAHBLTl
=
0
)
(
input
[
31
:
0
]
CAHBLTOI,
input
CAHBLTII,
output
wire
[
16
:
0
]
CAHBLTlI,
output
wire
[
15
:
0
]
CAHBLTOl,
output
wire
[
31
:
0
]
CAHBLTIl,
output
wire
CAHBLTll
)
;
localparam
CAHBLTO0
=
16
'b
0000000000000001
;
localparam
CAHBLTI0
=
16
'b
0000000000000010
;
localparam
CAHBLTl0
=
16
'b
0000000000000100
;
localparam
CAHBLTO1
=
16
'b
0000000000001000
;
localparam
CAHBLTI1
=
16
'b
0000000000010000
;
localparam
CAHBLTl1
=
16
'b
0000000000100000
;
localparam
CAHBLTOOI
=
16
'b
0000000001000000
;
localparam
CAHBLTIOI
=
16
'b
0000000010000000
;
localparam
CAHBLTlOI
=
16
'b
0000000100000000
;
localparam
CAHBLTOII
=
16
'b
0000001000000000
;
localparam
CAHBLTIII
=
16
'b
0000010000000000
;
localparam
CAHBLTlII
=
16
'b
0000100000000000
;
localparam
CAHBLTOlI
=
16
'b
0001000000000000
;
localparam
CAHBLTIlI
=
16
'b
0010000000000000
;
localparam
CAHBLTllI
=
16
'b
0100000000000000
;
localparam
CAHBLTO0I
=
16
'b
1000000000000000
;
localparam
CAHBLTI0I
=
16
'b
0000000000000001
;
localparam
CAHBLTl0I
=
16
'b
0000000000000010
;
localparam
CAHBLTO1I
=
16
'b
0000000000000100
;
localparam
CAHBLTI1I
=
16
'b
0000000000001000
;
localparam
CAHBLTl1I
=
16
'b
0000000000010000
;
localparam
CAHBLTOOl
=
16
'b
0000000000100000
;
localparam
CAHBLTIOl
=
16
'b
0000000001000000
;
localparam
CAHBLTlOl
=
16
'b
0000000010000000
;
localparam
CAHBLTOIl
=
16
'b
0000000100000000
;
localparam
CAHBLTIIl
=
16
'b
0000001000000000
;
localparam
CAHBLTlIl
=
16
'b
0000010000000000
;
localparam
CAHBLTOll
=
16
'b
0000100000000000
;
localparam
CAHBLTIll
=
16
'b
0001000000000000
;
localparam
CAHBLTlll
=
16
'b
0010000000000000
;
localparam
CAHBLTO0l
=
16
'b
0100000000000000
;
localparam
CAHBLTI0l
=
16
'b
1000000000000000
;
localparam
CAHBLTl0l
=
16
'b
0000000000000000
;
generate
begin
:
CAHBLTO1l
genvar
CAHBLTI1l
,
CAHBLTl1l
;
reg
[
15
:
0
]
CAHBLTOO0
;
reg
[
15
:
0
]
CAHBLTIO0
;
reg
CAHBLTlO0
;
reg
[
31
:
0
]
CAHBLTOI0
;
wire
[
16
:
0
]
CAHBLTII0
;
if
(
MODE_CFG
==
0
)
begin
:
CAHBLTlI0
wire
[
3
:
0
]
CAHBLTOl0
;
assign
CAHBLTOl0
=
CAHBLTOI
[
31
:
28
]
;
always
@(*)
begin
CAHBLTOI0
[
31
:
0
]
=
CAHBLTOI
[
31
:
0
]
;
CAHBLTIO0
[
15
:
0
]
=
CAHBLTl0l
;
CAHBLTlO0
=
1
'b
0
;
case
(
CAHBLTOl0
)
4
'h
0
:
begin
if
(
CAHBLTII
==
1
'b
0
)
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO0
;
else
begin
CAHBLTOI0
[
28
]
=
1
'b
1
;
CAHBLTOO0
[
15
:
0
]
=
CAHBLTI0
;
end
end
4
'h
1
:
begin
if
(
CAHBLTII
==
1
'b
0
)
CAHBLTOO0
[
15
:
0
]
=
CAHBLTI0
;
else
begin
CAHBLTOI0
[
28
]
=
1
'b
0
;
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO0
;
end
end
4
'h
2
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTl0
;
4
'h
3
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO1
;
4
'h
4
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTI1
;
4
'h
5
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTl1
;
4
'h
6
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTOOI
;
4
'h
7
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTIOI
;
4
'h
8
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTlOI
;
4
'h
9
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTOII
;
4
'h
A
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTIII
;
4
'h
B
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTlII
;
4
'h
C
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTOlI
;
4
'h
D
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTIlI
;
4
'h
E
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTllI
;
4
'h
F
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO0I
;
endcase
end
assign
CAHBLTll
=
1
'b
0
;
end
else
if
(
MODE_CFG
==
1
)
begin
:
CAHBLTIl0
wire
[
3
:
0
]
CAHBLTll0
;
wire
CAHBLTO00
;
wire
CAHBLTI00
;
wire
[
3
:
0
]
CAHBLTl00
;
assign
CAHBLTO00
=
(
CAHBLTOI
[
31
]
==
1
'b
1
)
;
assign
CAHBLTI00
=
(
CAHBLTOI
[
30
:
20
]
==
11
'h
000
)
;
assign
CAHBLTll0
=
CAHBLTOI
[
19
:
16
]
;
assign
CAHBLTl00
=
CAHBLTOI
[
15
:
12
]
;
always
@(*)
begin
CAHBLTOI0
[
31
:
0
]
=
CAHBLTOI
[
31
:
0
]
;
CAHBLTlO0
=
1
'b
0
;
CAHBLTIO0
[
15
:
0
]
=
CAHBLTl0l
;
CAHBLTOO0
[
15
:
0
]
=
CAHBLTl0l
;
if
(
CAHBLTO00
)
begin
CAHBLTlO0
=
1
'b
1
;
end
else
if
(
CAHBLTI00
)
begin
case
(
CAHBLTll0
)
4
'h
0
:
begin
if
(
CAHBLTII
==
1
'b
0
)
begin
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO0
;
end
else
begin
CAHBLTOI0
[
16
]
=
1
'b
1
;
CAHBLTOO0
[
15
:
0
]
=
CAHBLTI0
;
end
end
4
'h
1
:
begin
if
(
CAHBLTII
==
1
'b
0
)
begin
CAHBLTOO0
[
15
:
0
]
=
CAHBLTI0
;
end
else
begin
CAHBLTOI0
[
16
]
=
1
'b
0
;
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO0
;
end
end
4
'h
2
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTl0
;
4
'h
3
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO1
;
4
'h
4
:
begin
case
(
CAHBLTl00
)
4
'h
0
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTI0I
;
4
'h
1
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTl0I
;
4
'h
2
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTO1I
;
4
'h
3
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTI1I
;
4
'h
4
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTl1I
;
4
'h
5
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTOOl
;
4
'h
6
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTIOl
;
4
'h
7
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTlOl
;
4
'h
8
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTOIl
;
4
'h
9
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTIIl
;
4
'h
a
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTlIl
;
4
'h
b
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTOll
;
4
'h
c
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTIll
;
4
'h
d
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTlll
;
4
'h
e
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTO0l
;
4
'h
f
:
CAHBLTIO0
[
15
:
0
]
=
CAHBLTI0l
;
endcase
end
4
'h
5
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTl1
;
4
'h
6
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTOOI
;
4
'h
7
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTIOI
;
4
'h
8
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTlOI
;
4
'h
9
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTOII
;
4
'h
a
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTIII
;
4
'h
b
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTlII
;
4
'h
c
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTOlI
;
4
'h
d
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTIlI
;
4
'h
e
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTllI
;
4
'h
f
:
CAHBLTOO0
[
15
:
0
]
=
CAHBLTO0I
;
endcase
end
end
assign
CAHBLTll
=
CAHBLTO00
==
1
'b
0
&
CAHBLTI00
==
1
'b
0
;
end
assign
CAHBLTII0
[
16
:
0
]
=
{
CAHBLTlO0
,
CAHBLTOO0
[
15
:
0
]
}
;
assign
CAHBLTIl
[
31
:
0
]
=
CAHBLTOI0
[
31
:
0
]
;
assign
CAHBLTlI
[
16
:
0
]
=
CAHBLTII0
[
16
:
0
]
;
assign
CAHBLTOl
=
CAHBLTIO0
[
15
:
0
]
;
end
endgenerate
endmodule
