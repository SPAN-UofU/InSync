// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 10Feb10		Production Release Version 3.1
// SVN Revision Information:
// SVN $Revision: 11955 $
// SVN $Date: 2010-01-30 15:35:13 -0800 (Sat, 30 Jan 2010) $
`timescale 1ns/1ps
module
CAHBLTllO0
#
(
parameter
[
0
:
0
]
MODE_CFG
=
0
,
parameter
[
15
:
0
]
CAHBLTO0O0
=
0
,
parameter
[
15
:
0
]
CAHBLTI0O0
=
0
)
(
input
HCLK,
input
HRESETN,
output
wire
CAHBLTO1Il,
input
[
15
:
0
]
CAHBLTl0O0,
input
[
15
:
0
]
CAHBLTO1O0,
input
[
1
:
0
]
CAHBLTOl1,
input
[
1
:
0
]
CAHBLTIOll,
input
[
1
:
0
]
CAHBLTlOll,
output
reg
[
1
:
0
]
CAHBLTOIll,
output
reg
[
1
:
0
]
CAHBLTIIll,
output
reg
[
1
:
0
]
CAHBLTlIll,
input
[
31
:
0
]
CAHBLTOlll,
input
CAHBLTll1,
input
[
2
:
0
]
CAHBLTIlll,
input
CAHBLTllll,
input
CAHBLTO0ll,
input
[
31
:
0
]
CAHBLTI0ll,
input
CAHBLTO01,
input
[
2
:
0
]
CAHBLTl0ll,
input
CAHBLTO1ll,
input
CAHBLTI1ll,
input
[
31
:
0
]
HWDATA_M0,
input
[
31
:
0
]
HWDATA_M1,
output
wire
[
15
:
0
]
CAHBLTll0l,
output
wire
[
15
:
0
]
CAHBLTO00l,
output
wire
[
11
:
0
]
CAHBLTI00l,
output
wire
[
31
:
0
]
CAHBLTl00l
)
;
localparam
[
4
:
0
]
CAHBLTI1O0
=
16
;
localparam
CAHBLTl1ll
=
1
'b
0
;
localparam
CAHBLTOlOI
=
2
'b
00
;
reg
[
15
:
0
]
CAHBLTl1O0
;
wire
[
CAHBLTI1O0
-
1
:
0
]
CAHBLTOOI0
;
reg
CAHBLTIOI0
;
reg
[
31
:
0
]
CAHBLTlOI0
;
reg
[
2
:
0
]
CAHBLTOII0
;
reg
CAHBLTIII0
;
reg
CAHBLTlII0
;
wire
[
1
:
0
]
CAHBLTOlI0
;
wire
CAHBLTIlI0
;
wire
CAHBLTOl1l
;
wire
[
1
:
0
]
CAHBLTOO0l
;
reg
[
1
:
0
]
CAHBLTIO0l
;
reg
CAHBLTlO0l
;
wire
CAHBLTOI0l
;
reg
CAHBLTII0l
;
wire
CAHBLTllI0
;
reg
[
31
:
0
]
CAHBLTO0I0
;
wire
[
15
:
0
]
CAHBLTI0I0
;
wire
[
15
:
0
]
CAHBLTl0I0
;
CAHBLTlI1
CAHBLTO1I0
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTOl1
(
CAHBLTOl1
)
,
.CAHBLTIl1
(
CAHBLTOl1l
)
,
.CAHBLTll1
(
CAHBLTll1
)
,
.CAHBLTO01
(
CAHBLTO01
)
,
.CAHBLTI01
(
CAHBLTOO0l
)
)
;
generate
begin
:
CAHBLTI1I0
genvar
CAHBLTl1I0
;
for
(
CAHBLTl1I0
=
0
;
CAHBLTl1I0
<
CAHBLTI1O0
;
CAHBLTl1I0
=
CAHBLTl1I0
+
1
)
begin
:
CAHBLTOOl0
if
(
CAHBLTO0O0
[
CAHBLTl1I0
]
==
0
)
begin
assign
CAHBLTI0I0
[
CAHBLTl1I0
]
=
1
'b
0
;
end
else
if
(
CAHBLTO0O0
[
CAHBLTl1I0
]
==
1
)
begin
assign
CAHBLTI0I0
[
CAHBLTl1I0
]
=
CAHBLTl0O0
[
CAHBLTl1I0
]
;
end
if
(
CAHBLTI0O0
[
CAHBLTl1I0
]
==
0
)
begin
assign
CAHBLTl0I0
[
CAHBLTl1I0
]
=
1
'b
0
;
end
else
if
(
CAHBLTI0O0
[
CAHBLTl1I0
]
==
1
)
begin
assign
CAHBLTl0I0
[
CAHBLTl1I0
]
=
CAHBLTO1O0
[
CAHBLTl1I0
]
;
end
end
end
endgenerate
always
@(*)
begin
casez
(
CAHBLTOO0l
)
2
'b
?1
:
begin
CAHBLTIOI0
=
1
'b
1
;
CAHBLTl1O0
=
CAHBLTI0I0
;
CAHBLTII0l
=
CAHBLTllll
;
CAHBLTOII0
=
CAHBLTIlll
;
CAHBLTIII0
=
CAHBLTO0ll
;
CAHBLTlOI0
=
CAHBLTOlll
;
CAHBLTlII0
=
CAHBLTll1
;
CAHBLTlO0l
=
CAHBLTlOll
[
0
]
;
end
2
'b
1?
:
begin
CAHBLTIOI0
=
1
'b
1
;
CAHBLTl1O0
=
CAHBLTl0I0
;
CAHBLTII0l
=
CAHBLTO1ll
;
CAHBLTOII0
=
CAHBLTl0ll
;
CAHBLTIII0
=
CAHBLTI1ll
;
CAHBLTlOI0
=
CAHBLTI0ll
;
CAHBLTlII0
=
CAHBLTO01
;
CAHBLTlO0l
=
CAHBLTlOll
[
1
]
;
end
default
:
begin
CAHBLTIOI0
=
1
'b
0
;
CAHBLTl1O0
=
16
'b
0
;
CAHBLTII0l
=
CAHBLTl1ll
;
CAHBLTOII0
=
3
'b
000
;
CAHBLTIII0
=
1
'b
0
;
CAHBLTlOI0
=
32
'h
0
;
CAHBLTlII0
=
1
'b
0
;
CAHBLTlO0l
=
1
'b
1
;
end
endcase
end
assign
CAHBLTOOI0
[
15
:
0
]
=
{
16
{
CAHBLTIOI0
}
}
&
CAHBLTl1O0
[
15
:
0
]
;
assign
CAHBLTOI0l
=
|
(
CAHBLTOO0l
&
CAHBLTIOll
)
;
assign
CAHBLTOlI0
[
1
]
=
CAHBLTII0l
&&
(
CAHBLTlO0l
||
CAHBLTOI0l
)
;
assign
CAHBLTIlI0
=
CAHBLTOl1l
;
assign
CAHBLTO1Il
=
CAHBLTOl1l
;
always
@
(
posedge
HCLK
or
negedge
HRESETN
)
begin
if
(
!
HRESETN
)
CAHBLTIO0l
<=
CAHBLTOlOI
;
else
if
(
CAHBLTIlI0
)
CAHBLTIO0l
<=
CAHBLTOO0l
;
end
always
@(*)
begin
casez
(
CAHBLTIO0l
)
2
'b
?1
:
begin
CAHBLTO0I0
=
HWDATA_M0
;
end
2
'b
1?
:
begin
CAHBLTO0I0
=
HWDATA_M1
;
end
default
:
begin
CAHBLTO0I0
=
32
'h
0
;
end
endcase
end
always
@(*)
begin
CAHBLTlIll
=
2
'b
00
;
casez
(
CAHBLTIO0l
)
2
'b
?1
:
begin
CAHBLTlIll
[
0
]
=
CAHBLTllI0
;
end
2
'b
1?
:
begin
CAHBLTlIll
[
1
]
=
CAHBLTllI0
;
end
default
:
begin
CAHBLTlIll
=
2
'b
00
;
end
endcase
end
always
@(*)
begin
if
(
CAHBLTOl1
[
0
]
&&
!
CAHBLTOO0l
[
0
]
)
CAHBLTOIll
[
0
]
=
1
'b
0
;
else
if
(
CAHBLTOl1
[
0
]
&&
CAHBLTOO0l
[
0
]
)
CAHBLTOIll
[
0
]
=
CAHBLTOl1l
;
else
CAHBLTOIll
[
0
]
=
1
'b
1
;
end
always
@(*)
begin
if
(
CAHBLTOl1
[
1
]
&&
!
CAHBLTOO0l
[
1
]
)
CAHBLTOIll
[
1
]
=
1
'b
0
;
else
if
(
CAHBLTOl1
[
1
]
&&
CAHBLTOO0l
[
1
]
)
CAHBLTOIll
[
1
]
=
CAHBLTOl1l
;
else
CAHBLTOIll
[
1
]
=
1
'b
1
;
end
always
@(*)
begin
if
(
CAHBLTIOll
[
0
]
&&
!
CAHBLTIO0l
[
0
]
)
CAHBLTIIll
[
0
]
=
1
'b
0
;
else
if
(
CAHBLTIOll
[
0
]
&&
CAHBLTIO0l
[
0
]
)
CAHBLTIIll
[
0
]
=
CAHBLTOl1l
;
else
CAHBLTIIll
[
0
]
=
1
'b
1
;
end
always
@(*)
begin
if
(
CAHBLTIOll
[
1
]
&&
!
CAHBLTIO0l
[
1
]
)
CAHBLTIIll
[
1
]
=
1
'b
0
;
else
if
(
CAHBLTIOll
[
1
]
&&
CAHBLTIO0l
[
1
]
)
CAHBLTIIll
[
1
]
=
CAHBLTOl1l
;
else
CAHBLTIIll
[
1
]
=
1
'b
1
;
end
assign
CAHBLTOlI0
[
0
]
=
1
'b
0
;
CAHBLTOl0l
#
(
.MODE_CFG
(
MODE_CFG
)
)
CAHBLTIOl0
(
.HCLK
(
HCLK
)
,
.HRESETN
(
HRESETN
)
,
.CAHBLTI0OI
(
CAHBLTlOI0
)
,
.CAHBLTI1Il
(
CAHBLTOOI0
)
,
.CAHBLTO1OI
(
CAHBLTOII0
)
,
.CAHBLTIl0l
(
CAHBLTIlI0
)
,
.CAHBLTI1OI
(
CAHBLTOlI0
)
,
.CAHBLTl1OI
(
CAHBLTIII0
)
,
.CAHBLTl1Il
(
CAHBLTO0I0
)
,
.CAHBLTIOII
(
)
,
.CAHBLTOOII
(
CAHBLTllI0
)
,
.CAHBLTO1Il
(
CAHBLTOl1l
)
,
.CAHBLTll0l
(
CAHBLTll0l
)
,
.CAHBLTO00l
(
CAHBLTO00l
)
,
.CAHBLTI00l
(
CAHBLTI00l
)
,
.CAHBLTl00l
(
CAHBLTl00l
)
)
;
endmodule
